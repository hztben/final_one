��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8F�:9 R�ibD�鶗9�1_>Y���4$MX:T7�q��N=����w�XEE���?��&��i��(��c}��&��>aӭt��fw�5)���; ��H����Do�6	��gy]њs���Bm��.�E�e��Ļ�60��NP��ب��Wx�z��Ir$%;M�I�Z�<6b|��m��P?�0<s��w/�8J0���:��T��I�;<�l�Yy\�7Y(
�����I�u�� ,uQY��j	����6	I��4�H���[�0;�F�$�ȣ�3�+�6!�u��׬�2~���4�kWf�2��]o�*��L#��z��'ى�.E��|��s�P<,i�a]���J����~TVhӑ�l�s&������DT�ND�5q�gl	�7C��r9��x�o�cy��:���w2�&�y�`�"�����W�+�;��g\�h���Ȫ�T��9{�E�#T�y0�S�LC�ۆ���k$;���9K�Q0��� ���Ɩ�o��|4����[�K���T)0�W�����������mh ���#xh�SH�]^e�M�Ǚfmv�~��0���6� ����З�55�Ac�N�P- ���uN��1sLcb���
T�~�\�Y�4��&'�%R6hP���A5��$���N���If�3wz��?b��Q4_��)7��x����'�C�9��~�w��<��qzcA��앣#�9Ö������ń�J�OQ��Z��8����29K��"/������F�[����	6>�kg��ߞ��]HV�pG�y��	��g�G�j]�e���:�M�o��%I���T���+N2A�H?h1|�U�{�ah�V���¬�k҇�E|����r��(^�ȱ�d@"��j��S�m9��3�e��uˎ�1d��kC �)�S�	B<��fΐd��<�e��L�����t;#�z{�Z��>�w��hA��|�)�b�j>��px�)a�����a�>j&��$�Q~W�|��e1�?�nd!TO��b�Q���Y�{�)���	�e�kP�j(}�(g$n:��e
��o�O:���5�p�쏦N|&��2��Lm��y�M���/����h�|��a��B��L��GI_�G������HÅ��_�q�_��*w��"(2�}P�oU{D�k���~ßC���ܻ�*{��<��/�2z��H�6���z�?����z��o,'����a_C����̙��d�v�%�����ɝ�.O�^���?�͜��g/�JY�D2�H���i�I�Vb�b�]��ZY;%�L����a�VzQ�nz�m���Y6J�\����$Z�9��y�9,�ո��KzrU��#k��J D�6�MP	~2���5�y��L���H�1�Xy�Q7�Yn�2����Ô�1���:�y&�ݗ�z���i-�H1�X�{����DkU��0^`1ֻ4��[.D���J����`�J|6���2�.��A�1ս��yM<�L���ߓ�hdw�����rΉ~Q���!�_o�Av�Kp2�s+���Ԥk2d��Wq�:%um#����Mb��T;Q�x�W{ܗ[�1�e_녛���W�*��	-�>���c<��+9(��}�=����L��	�<B��8S��.B�	:�bH6�;��I�b��h ;
[K���OH�"��_ �d5���=��d�}qmc�����\��9����E��"���wU���>���܄G_��-��Z��%,�7b�!��ejU�{�r��н*�pS2f�L��|���v�!Ri�=��_�������[ۇE�
5v��8�M���ǠKY�2TFX�e���j9��́DN��1�����n�D��x�i�v�;�U����!�k��b������6d)E-����O���K}
'`:cӕ!�rȄ��l!
�LX�3��H'j/q�(���W^��V!��^Zv��`�~��,7ߕE�4?4�	^�_�җ�t��P=�x˪��!I<�D�T�����F�s�_ �z^�ן�0�Û�Y�����S+�+N�Pa��S� �FU�%��5��a��xi�ҶaQ�n���z��D	��'��(�&pQ�(-���C�2�BÜW���޼��͕9�c�e?�M��]�����DI�X�._d��2���yyG=)�l�Y�ZD5'I�4,[��0S_��q}b�����q�0��nW&2��ۤӨ���E���ַ߈���(��@��@^F���E\�`=/�7ǫ��D�-ce�;P傿�a�#0�ev��lC�Ӫc�G��ʎ�)d���|����#���	޽��)��K��0� R'����'��lDϓ� �s���i��h���Ko����b;A�A�E�D���Wk�v�ɼ�ɶryc�����Zy������1�v����8����@E�r�nӬk֒����x����ǛD��s�Ө:���_Oi���������8f��=�p��G��� ��JFƋ�XQ���,�7�D����?�i�-�@RЅ����X}�Wmk�fp^���ߺ��t�(V�c���HK��]39����)t�1�t�c+����;�W|nt�'����:��{�J\G-��!�����/��B>�!|��mf�<����l#t�lyҬ_{O�vH�����CU~�i(�0��d��*��	��}^p0S�)�+��X`<�	E⑰�5u�^���@�z~�C�SG�p:�&��Ν�em\[sФ}��7�9*�$���05�I�Cĵ���7��>i/����	^v��ꙝ�*s��J��l�	�މ��vɖl�^�1f6+���+DQM����'���?×i���D.M`���ݑP��Oh�	ea��0�2��o~������P#�Zv��e��f��-�8bj ׀�V��ZJ)�)~��Vo�ޓ�ID�wʈx{W�?r�a�&����2^�K��������BS��@�_!�,�۹!�>_�X�Ø�48���V�L��c5Y��-�����A���w��z~� ���@�;c�0�IĮ����[_�oX I+%L�B2L�vp�/��c�жLX��k]�gsI��^l�^	8�@_��ו�,���(�H&�j|���5)�vL>�dÌu�{6��#�ߜvj��+_��ӗҒ���!">V���Z�������cX���f<#�&is�,Cu�=���%������ʍ{����f�v�hޘ֢�~�GΦF�@�i{C��om^�#)'$���sǴ-K�c��?#�#�x�H2���_�«H�C_5\�C!���DF�p����#W_qA��FU/�@�f�����C(�>銉�����E��I(�/e���bU��W�GEDKde��ǲ��!W��R��F�������t�w�X-�kMX}�6��G~����OE���H�<&��{H��L�����f;�l󭧵'�]�`��|���Ḋ�{�nq�u��a'䦥�$x}�'gϔ�fיx�q8��כ���M���y���Ϋ��՜T�cP���4�3�P�s������[-0hxK�q����ȍ��va��%ޠj��7�F�Z��gBo��t��\��3
�^�B$K9;#�	x�!ČEu.w�D��h���S�$ʎ T�^U��"���5 E�7�hi�����~�˽~�ZnMŽ��{�	�p�~�/W��kU#�~z�H�LMr���
���=��	qA�s�&S�����V7��s �D���i��6��%���g8P;ʗ��B�S�0xu��=���B�#��P��g��1�T���ޔ�o��X���$��c��I���� s�'�i�=ܲ���>R_�!�d�.?s�PJ�^��ˑ'�T}Z�nF�|�¼���޽�#��-����z��~�s�C����b�I ଀����L��_6p�+����\���{�x�x�>��'��@ *�6c�\>m�Y�g��Pqk  �@3���00�Sp�8�#e/�yc�������<l�R��\
>��J_����sZW����A�3����Z�Py?}�VM.���1<��kݑ��ؔ�@�����V���`��C\BPK�d�:)���X:;� %{HW��LJ��Ύ(��U3��]��~۷s���� �v���C�[�����#'.ƃ��e�ϡ$���?em����Q8�٘{t��ts5[C�Tfe')��Շ�M�U�H��5��?f��8R�t�AyٕEN����o�0�nf���_��H�ѭha뭞�:Z2+Z=T����
���c����DE�F�N��T�m՝X�C�Lyҽʷ������U�eT��/ׂ�b`d��^,�_�/
lD���%Q��%��tDQ��d��<�����Ut--h>�?�
!�Nv�p*3���ċǽ	�M(�qVeP�\�zI�rh��֣@{9h���T��L�=Q2��ou����y�
�o�S�2�8��#��=].1dL�g��Kτ��d?ɦ�I+y����}��9�,�t	�(�U�B���4��T�������{T�g�,���~��N���<����~x@���|{%x����7L��j�<P�'d�ޝ�H�%�ZD���������AN��ҘP������Xt1y.�sd���T���.V�c4E�U\�ľ�t�t�)~�YL�̽��"4^A5�D�3��ۏv�L�a���At�3=L��Ն��}���zĚL[38R"�|^���?�TA���td��+<�)ɖї��LR|ё�!v=��A_���~��z�%mxޫɷu��a�XJ$ҋ}5�J��}����z�һ�uV-kIr�a0�l��NjR{�y�^��UY$G�N�����$s��
(�Ý���N@!�o7+����$��M�Zo��T/����%E@'�߾�{����g�ypB�G�f�Z����3�vMoE������t���!��}�x"��}�c�<Rz%u74�L�e+�W���5A��g��VL�)���0d����E.�UPEP�
׬�pgwش�ZKU��Ko���?��F�������㪨���yT�ď��5@�8��#�`��	���S���so��
	�6g>/�nN����(i��>�F��h��x��?*ΈL�	Zaڿ��η��W;�QW�=m�G7qq�/q�HO�}��>��Y���=r>��aG���s#U�/�|?��N���.%?�#��iV�D��k��i$f�$%.8��SX]�!{y��r�r��ڕ7���a���s��Yb\DP�9d�o���� �����}�R�'��U�箱�C�"�4%!$�ܶ@~�=���}H�*]̥^pf𨯙�BS�X��	�b,k�}�ߵ��8qM�ʒ�2�WU�����IHGv��`4���r�~��ޮ/�KF�J���U=�Q#L�zLĥ���� �r��Q��x{o�ʥ0�6��:��^#Dz��f�����J�;�-y�&4�J�~ˈ'�)�I�������گ��C�=�-����NFP��5(`PJU�J��10�
��A�y��.�t�,���@7�� g��B��Næ���dc�@&b�6��^w�-�p>��Y
�cտa[�L�9Ns3l7Y�Z,��r�H��j2c���%�Bܚs�n�a�H�ϴP�C��)�>i!S�
���k��7Y3l��R/��d\rZu1 ����vo\���[?������%sG9݆�	&�8��2�/�t'7  H���!��5a��>�2;j�	dq�aO����^6��P�����.$~�;��S��!��@Se痩1ƟI��9���B�T� �ǐJC�CD;6*��*����F�L�����t�>v&h�J�����E
��%��d���ZdԌAϧ�<gh�M4}T_���{bn�s8���r�|�� �1;�R]�}#\{c>�^o��؉�®*�e_8lI�	��]P$U�q^	�0g-^�O�K������R�� K�I��_3-T�I[V�8h}�P5��%�rҍ�+��,����g�/A{�� �������*&�<����o[%G�F�Ҍb�91#.��"a��A;�ʣ=���Fva=bM�~E��81J,$���9$���J=���o���g�2( ~O�[�M�a(�-���\80GǞ]��ҹ�ϒI�	���d����F3ˏ�F2�C��+�'&F�i�����~�w�R^J�P�9����P���"��ٛ��~JC�I(S߯h�˜R�J�R0��V�C���)W���������Tq<r.��L���b�wdtH�_.��pm[`:[sngu���mn�$h�A��h��<��m9�Eɽ3h���M�l�|�W����v�M6]��g�nr��߁͑�V/�=���9��1�`X����:{J��fvT�JNR��#�8����Ѹ�
c�w	s���C�g��;�F뀬o~�)W(=cD���$)�Y���0xa��wA8�^P7_�Ge��4��}m��/-�R�R�WL:.���9��!��@)��!b�L]!���������5�p�D����3�'x�a������L��H&|���*��a\
�ҊU���Xjp񽵽��3MN�V�ȫ�.��ۢ�k|ϲ�Z�3J��C��ܾ�sX��_A���ݡ��(�R}�ե
�f?��M>�ag	�� ��Hv�>`��:>��J�\V�E\�����5��W���H��łt����AID���x	�B[�K���	�BK����;�U 'o\�ǅ*�=�Rz+� �0O�d�0�u���jEK��w�S^\_���H���hC-q��G��?�7i���a'�2$D2z�,R�0���1��7�'_����	��:�|�N����Y��b�ue��g�$Ω1\ݱ8/�����f�jw��ɴ�`Z��M�'�l� Ϸ����	�	�3�1x�����e�Z���:/��s��.�5�_�x�,.t% ~�p�p�r�3N�sĵ�c!%�7I�R�����	l�|
�@����� �i�˶#ɍ�S�jG'�]�Wn�ðLj��>��#�j�ǖ�J\���!���m=���ݙ7ǀR_�ٛe�{�i��1X|g�Ud�Z�*��-��Z�}*%��©���z��܈9a��u�̻	�)����&�<>�ڷ�����駚t��"�ᑹ�]���Ŷ\���`�/^pf+Y�]��<g����eO3���[���F�<v�ߵ#O���<���:©Oi2�%6�(��jzC��&+�(�'P蓫��j��5uqc�������/m�Gh��G�d1OB���/!d�g�vkw�4���G>��&�C��,g�A��0Z6V�h޵���0��H�ѐ�a2l��#�HC%)�
GU�z�-��iq��ՆD���V
����c��ޮ��9\6��^��YE^ȃq�G/0����Md(@��#�5AE���-ӓ����c�^Ho��C��{�]G�$)�d��;
o��;�!�4��G`L$��v<����"V�������
��I�2I���q��#1����A���(,�m�)Z˭ڝ��]>��_s�.t\- ���"��VrBwZ ��!��Wzѫ�Y8�]��a�z_��h��7yt�����c8 �[W(�w	���W �Qt�(`q�i<	I�Z�d>�*�O�h�����"nX��g���,�����Z*2;ã�E�5ܴ���bb�_�AX�_w��iI�=��L�=]����&��a�Y�(Z�Y)H7Z��Ths���$����-�̷��W$�v6R�!i��!1���Y���/�E����dfVJ�1�Ö����y��q��o�|ԋ�pw,���᱒��j��j�j�.0���z�?�!��y!:��@sG'�F!�E�r%�YE?Sdf�R�^����w�,��b�:����04Υ�!
.5���f�����	<�'�ݾ�*����~����b4�^jY��ΧgoC��(,����]��.��8�g��г-������� ��ѧ��7��D�s;�����F�/�P]P|��zX�@�V��3�����4�*+(��\�M5�kJ�A1�-RR��.�Ta�R{��m�H���w�³��E��PT��6�D
��zP���`�;#3�б�R�E�pԒө(5]�������EJ��v4~X�#OC҅����j�XܕBڬ0?&�ʽ��@[m[:�t
�w����V�	�f5۪xI�w�T���S�R'�}Ux�"c��̨2^k�[砅��p��R�|m	�@C6���F�)A@�.@��|rH�(�f\�q�E�s�t�δo�����qL�H��{�K)�3�t�W� �o+?�#��m��+�%����߉T-<�t�L�RɪA��L#�$O(r<KF-�
Ǡ�$b?��c|w��R��i���wM����Ǫ�<�l�+��d,,�AX�a�D˟�NK!�n�f-t�W��}�1.ڿ��NiK^0�sh3��(q���&����Nʸ.m���m=���}���ڒy���8*k>��櫡�l�69�c�[^h�5ׁ&nv�Tr���|�u�k���j���H��.f��k4ü!K��@F�C�7?�zW	�LIOT�P*n.2��L9�(~���ђv��k�A6�[���
�ty��k���ʪwp$�n���˷W,C�۪�����/o2�rR��>N�w��񠼭�'GV�o����3�dޠ�һE���hP��ޜ�e ����]x1n���I�)�p^I�ؐ��������G���칅Ȯܖ��DA�4z�OK��2(�I`�\�c��-��йぞ4
j�`��ϛ�]����2-����i�[%5y����bu�nK�*ԆÃsu{���w��2�58�bzmǒ?(�{�6m5*&>�����E�W�6Zra���#%��Q
�lS�%��h."��Ix���@a(�q�'"75-x��Ч^��V?i�9�X��5����kcM�R{43��Ʊ���J�����hɝ�J��t.d�tP�K�=ђ0�)ȱ��%R�!�S y���޶�i�1dIb�����1�/�e'!Oh�=�4�F�+�+��v�����1@9�✼	��e��,1�PЂ�^�)��2��[����%W�yp�9�[�n������N"�S�l�_#>G	my�Jp5-�%��@�/O<����9��1�㳂�AJ�$'���䶫��̀4�|<c���X7:u}���	� J���$g�,)��E�j<ˇAx[���\	��1"]��e��E��Xv�Mo ��$v��P	�`Ŗ�I��L��z��~�]$�S�G�ڐN���$s��Y�ɬ������|OS�%���/$��?�d��ְ�&ʿ�P�D/r�r(���z�O��	_@��nmjGW�q.�f��I��5��M�B�ym�l�I�U�I�i������yPt頖�e�Y�TD���K�4L���'r�mk�E�����$��kDSԢ�4�2�kբ;���r���#�|��ԁ".�9�9w�Bm�]��J�?L��6٧��p6�r��vݷ����nĨ�nYdB�Q?r\7~�si��j��t!��n��>�ç@��Lb�ysOr�����A�p�/ƃ|X�/���p�H��7*�rո�@��~v�a)h��ƞS�&�9�����QI�@6�Ns��itKM�n���k���ɑլ������)s�k	���v��3�]zJ-��X��K��N2�VC�o����I���9+��k���d.�������w+��{i�*2�Ŝ��e�`9OE�0Z�f�-�����˥�:˛c���B����Ǎx)�w;7�'<�m�ax+�'kD��]�i�� �u�%��	s���C/�G�Џ[pG����=��!�uFT9�7g��O��h��0�o*�y���F��~���}���⥪�sp���r�<��"����pK����}o1莃��*�w/� ���m�3d�eߓr��" f�D�0/v�r��r]ꐰC~�~��lG2"��b02M+xQK3e[������ӪC��H_���A��l?#Q�&א�ŵ�2YH���Q4sv3Gڒ���D�B�Y��G.�q/��B��1#��K�-�s�ߡ��<���ɋ?L�r�KI�9�{�}y�D�ѕ�I�
2{<�k&�6�W�:a�QOƉb��7O�0�!�r�g(�d��&�\�J��WEh|�,[KF0b|�k4���op���+����JJS"�0��44���]K��T��ݜ�/g� br_��LU��>�!����(�s���*;[QM��x�$�n,��1u�Α�d�<%VyV.bN�e�n/LӅ՚-���/Fh.Z(��nc�(/�Jg��!�-Ľ�y9�)<a��a��E�}�Q׼ўT�h�@}�bKaQLs~ʺ6#���w�t���y��V�I�ջ]��r�{Y��?���ɉ�RV�\���˛t=P� ���/���Z�y�m�d+4��ӷhDڪ�K���2���𖑭 ��qbӊn�F ���9(�l���~�}93g�� %|��}PZ�V�6�ˋ��PT\�����g�d����(�w�r�յ?^��[꟬��[æ��L�JLV�9(��|GyNyWҺ�r�UE��OF�C��J�K�;Fq��1�XS��E��f,��%BpX}�V�����`�X6!�A�� �G/�Ġg6<�kGv��v��x�M�$U�gSQKAm��OZr �_�$��$g6t�JͶ&���-.��-��_[��]L��;��Yk�hgsm�-@��Q�Xo� o�E�\��G�ddֿ�}�vB�N��O���[]T�������!Q�LN��G��l��1QI�f�}��K��u,��U�͠O}'C�I��l$�� 3�W'���Z�~�j��Bab�:�L����Ց��P�b��+ ��'`flWpx�������tR��40�I�����zZ�.Xu\&���)�� ��\����`���0*�h�aᢌj�!�^�~{��{􃿼��՘*�6qI��к�J0�n��b��Ô<%�֌d�4g��*0�.���|ѝol�$���a��/�5E)c��������z�WL ��S>'�bm�a��F�q4��T�'��h+j[q!d^��Z͒g��2e���|�Q/�/�_���������yt�'��B?"\���%k+?p�Q>`�P����Q������3��o���U�ua��Ş�_R�H�(c���TP#�	�е��5z��T�`��U���$�Y�{Ф���17F��/5�����2O�,�JgΝb����D�%[vPQ��Y�i�����/��V���=�7I�x�\0�g�;&W}�m�`Vs�{��-^��L��R�*����>��7U�4i���#��«7����H�/��ݫ�><-]���[�*�)Ҵ��<a/yl��g
��4*I�3����s�0��춏�O���F�&y;����$*)��Pe~i�F#��۬f����'{h�MS.y�1U..��cB��Y�W�2��5��u؟ٳBpR�Y�L)j0G�%g,���[/D{�kD5�����J�O�7ڷ!l�&tܢ-ͫD�����6�vb�t3*@uV[�ى�vB�)J���䎷Uf�R�H��|]`SX@��q��*5�q��"ٸ���.c4[���"1:<X���>�D&E2���)��e�B�< ~�A�St��3z.)�e�!=��+��B�/�Q�4
��񝋃MR�b�tgA{a���j�C�L���NJ��o ���ɐ�W]�^�.�0����Y��ٿ�@UP5�MV7��
"��>'sr�qۚ_��A}� ���z�|r��+HR�N5�2c̓H+/�0��,����f.�ٮ���� `9���y���B@�!D�����j�鄦���w��ç�){>+�W޲�q�P��񼯡a�'KV�6���C�:Ϡ�O| a�L�����a���hg���ڔ#���➳7 �O�	f]�QJ��J4����)P"pL.?��e�>ܫq_����E��2�s^؀d�:~";cj���CAEz�q�nPm� ��~��h�+{���;�p�n�ϫ�we4�S��Z ��JF#�D�.W�s���΅�	n���v*:/�2�"�O�|�H�f �!4*C	��I=�tF�a^�-H��	�wc���7�����^�N`�Lh�B�l��O�Þ}o�_���V�#��E2���l�
�=�O��۟�>r�JRT��v+���牟�DB9|\���&�[��$����n���;?���Éh	��Q�J_�弩��^7X��}v�rMj_�����=n�3f����IZ�+�[��G�a�H&|FT����4g]7*0Q2�;�V�{Z8����������B�;L�@^�$z����a�����x	2�Q���ܪc*�rp��R7�>��{H�F�}M��i�$4�ߗ������q=Y�J��� ����$�o�
�q[	� yV�i�b+k@H�ʝ��C>�3��O0�K��"m�P-n��E�*{�u,�1~�U�pK�j�5^1Դ��ńA;��6�w�L�O\�i�nh�'5:/���x��25+Wo֑�Eb<{23H��bG|���r_�hfh�|9���e�A8��F�	����n�����AsyI��H������ӆk�ޅt�!�}�dL���yD�3������H2c�H�?�������(�u��!@v�@^r��P�w��S�Z.i��q�l�c��uȬ|��.��-��al����U�����?h4�0���<����ɽ��ml���4�KRG��\�V�u����E�@�].��cK��O�~��{Va���)�����k���R��rj�d��� a��l�<W�j1aH1X�h�vL�h�H�#� ��̛�*���4�k�츾۞7��.h�Ζ4�*Vf{O3���׷$s��`L���nӟ����7#��)���FW��u@`W�K�����и���0�K��j	�w�{�b�ַϭQ���3�H�A��,��S��h-ۣ��e:�E���q(P��ƈ�
X.��2dx`a�G�
�>�f?%h�X{]fX�&|��3�E#�]�2���Ъ*��7�Y�$Z|��U�iD��&M������٢g�G��¨2"q�����;LȄ��]Ш�qdT2Q������P���L,��r%�J����(G�[�_9s�	�Q]����t��_DO_"N�A&��_�U�(yu�8�L�&p��6>�D�>��N�ӿ�O���N̬9��x	�ܴe�U3���@��-���!U�rer�Q ]�4�N�%{k�#�$v���f�_��������H�Yb�.T��&e͍y�s���U4��]
����"逞N���V�#�J�Ӯ�#�]Tx1�)�JQ+0i���cO�1�͍�g��A��P���JB����w��k�����P�C�.9ө�����Ki3)�*k�@T��f��N�E��P_m]�i'��Vxɿ���9���R��A���e0A�@)�O�F�kCe=Q���G�`]�5Q��Z�䯂:��Q��|35���ܕ�q_u4�\��� U�Ο�Ȯ�6�G"7�#VA�+�������y� �Eo�k�>�����U񚐀��Ւ��#��]�������A�^�dz�O����_��!����[l�Z�m�tB�;b�U�M
���?���ȼ��XJڦ�N��t ��P!zJ!R�Av ^����ICM� ȏ�W���� t�,^�T��|�����6 �e͖3��r�r�F�iG3[G�]�Hf-�~*��J*��?3`Y<I�I��5�!�m{&�|3�{T+����m]���^$A�i<$�Qm)q�ڈ�KA�#=������O<ڻ�O@��,40$��Jw`�{f�59"�ӎt��)c:��k]Pb,p�Ʃ������o�C����k.R�"	�/�{V��w#�Zh	\����Hh����.ZK��	������W�{@��aPr�<��8Н�^⑃	d'�u;)�趣�Zܨ���-~@�:d�����|C'�a��x����yF^6����"��`��Q�\���9X�q�N�/L2���)X=ӨV;���H��~e�/��]��I�J�g=姯�����Ʊ�p�����n�l��1���ꡜ)���%a!� �R�Й��K��xIv#���}Upc�n|���S�$4:V�H`�X㒋���Gˆ}���,�Obv20q&�ڴ�s�ふU`�� "�Z�����F1��CC����g�n�<��#�lD|��D�A����,�#�؀�x�JC8r@�P��tZ�����i�m���f=�$k���~��a�䭡X����'�RI�V����M�Fry�Hd����tBO���P�3K��,x��{�9cm��ݎ0Jk
:Tz��}�M�߯{J�~>�Wڳ.�ǉ�wz�E���0s��^<.�;�(���%P�L%{}�'J�~$�:�hQ��`��7�Kz=�Ӑ�2�z�N8w)�cV ���E�q
2&)(�Y�e�ސ��qC��[;���i[�'N*W`�5�Q���r�Б���1|��r%�n'ɣ�b��7�e�7�K�L�+�|�X�4�� �\1�/�E�g{v�"(XY�o����ǈ��U��
�0���j�"���#�h[��o����B�T��U7��o��4��l;B�$u�3il7-�NC.�K�~p,6���/�0;BF3\�A84"V���l��.�n��DVyݗ��I���o^ߕNSM9�l����C�m�o��!+M�hW�n�~�)3G��ti�I�"Q�)������n��I��9�����S?�
��Lv����g���-y�#��7$�s��'�� ��+"Lݰd>o<b�\{5�7K��	(�d*��U�C�9�)+�o��iw.%����*��!��ޯ8Cӟv�7ld�?�H�4�S6'&շ�G��D�������N��ȞյR�I��U�%�쌚��aC���������F����iie��1��Pel���u����ZNAlE�_�Ï�V���Q8c�s�b</v>v,�¼ X݂��pώ!�`aԭ���X�¶�����ޤ�T*��k������Ő���&_1�(��: N�Oݲ��q+z�zz<��d4]{Caщ�ؒ�΃�毁�rB	{k�N���##�P�V�0�G2�[n���u�P�'m�z�O �t���'f�/�� �tj�M#�ߌ
p��7u3ӽ���RX.=�~�{�G��5۽!ȵ_c�p�>��u'X���#k��?�QfdRȭ��2�=�E�Y�	����S^� �U`*\��Jc���z��B�}V��Zk���m.o�se������UV�"���"�����hL/�0�|��g+7	;q�u�V�Pƛ�����ǡ-�ײ��w�\=�Bg�0��0Y�bWr
ӈ���!
��AX*e<c���|��.�4L �76<�jޑl#�0j�w�V�F��+&�&�����s�$��lMPb*q��0/�W��e�`1�y�2�}�V�ۄ\L���fꢹ��	��Ex���������rA+*����,�����&��IW��&���G��J�:";;�<���0e6�]o��;<Q `2�-�vSᾢ�f�{�R�`�t)��岫�J`,�������`��@m�Q�k�g�`�"\VC=�c��[����p[j `�0��[@��z���͎�H��;	�Ω�/�<\�օB�1A{�����Q̿��q?��`��L3�e�ֱ�+?:�r�|�{.I��J��IT�
v߳�˥wۍ�f�/mR8���ԓ�OA��B)֡S�nʾML�qW#���XO`g�Rr�T8M����� "ʀ�&��$E�RH�O�ɓ�	}�r���Ӆa�Ord������.�D)�R���9��e��=���18���;Jt�f���d�/NT��M6�]큟 �5�	�r���UyĎ6�������wX���
���k�)��U��v�
Ð�A#.�\�N"��X*?������K�n~;HN;o���ܭ��K5��$0MjC��y��U�q!��0y3�z�����:��%���������U:D��e6G\�6�x|��̱�
����������5���"77ƪ���S�D
]\_�P|Æ�(���7��oҊO1u,v��QbxT�̢�,�B�AK��a?�
!l	���Q��V���n��%�F�E��_�V��/lY�ri�~�PwI
�	���t�(��X8�~_վ�͇�K���W_�l�Ѐ?j�W��A<��3�,o�Y>�U��*v5x]�Ս��ʤ�h��H�����$�.�u>8�����QJ�2��Sl�'����F�A�
#�_8.��W��#Y戃��3�EaO�_Y��*�c��T��$�h�ǐ��\��j���s����%p¢_�]��&9��i��� q )�{�������]�I��
]Q�Bi�<4}�Э倴+�;=;tu�tf�*�-Y�̥%��9�.-�Mv��?�V:� r|D��z�����e.��zL��Ӻ���Q"J��4�1����*n��'�k�N�Tc04{���J/(ՋS.`�b!9�w�aG�¾%h�)
�N�{��F��R�.��i����*/�;���sZ5��1;��@vB7U#�ujGz�6�4�y�Bd@R�Y �(��a�j�"�&n�i��)3q��T��P������sV�4��D?�K���r�Y�[PA�%D�>�*3��uz��[<�濒=tQ�7$�c&V�zc*�p*�g���P/8Q��"��d������2��cΓ�v�_�}�c����sr�`V�{��c5��Yb�p",&8-�;1�Z�7��T��GS�+/��8>ۊ��s6�y���*U�Y���E�`ɷ7!{���I
e����8��D]Fģ�Xt����c�n��gXd@�J�u4�?8fy4�E|-��oh���n�<��dc�n����'�S�Ŵ��57�V|�o�B��HbDL�9�D�Ѐ,.����%M�� S�͸��=6^�xo�����/=˗�ό/�g��m���۹�E]���٧M��	|�G��l��5"�[����E
�^�|�,�]E���O�Fw>�|T;���|����.c��I���n�ق���z�K�X�Zc.Ѭd�,��vp�0�hh��T,2��v��v��vI�}MjW��0_�����O�Ny���m���K*��(�U ׂ��b�:2��a�t�.��X4�p=R��]N |$[Ŕ?�!�o-`U�-Ҥ�G��'<����፻�.9�"�����e��	b,��K�h��mX�N��� {E>JﻉK�	���w҃#�]��48�!f�_~)Tw+�nZ�A8Jr���Ɖ�W	Ӡ�P����$���LAh�3K��/X���d'�N{�I���e5dm��@��	\�na���5�A�\ڎ���"q�-�f���9=o����.���`���F��d�#R�Xkp�����N폁�sD�wn0���xWаJ�Ѧ�`��=�9qC��Q�c�'�� ����J9!��*u)M���I�n��|��Mx+)������i�$�}]ہf�x������Ź�xc�'��I����՝G���(�W)���L�V,�jt@�a`�_|�z���� ���i P'��}���5�e�6'��a�)�,}��'$1f����/�N�k3�鄲���n����P��d�}��OMa#'����s{���LQ	�3`e?�g��;_�Ͷe&�y�`�g/����.�J�-U|Y̫��Y�r��f�3�Nr"�	��㍗��w���ɬ���=��`��|���U �i��f!�aA�°d<�%6p���"Aӫ�}�~:'|����0�{�}+	�Ru͟/����Nh�3�3�[��d�uc`����	���PR�� _�C���%~rgU[�CR^DBq��U/i񉢄?^��;����A߂"�N'#6��Cyo@�<��QTWW����!]��ϝ����X皾<j�dz�'ˉ�0"є�gX��G}�ه46:�Ā���ɝ�m���X�C,y/۬�1�%��nY�a(��	�A�<��2�dͼ�"zꈝpG�NE� � C��(U����m�U���M.ҵ���,��Bc��Bw���[�=�������y#�+�l�Ӽ8���471/�՚�z�H��̚'h&�~��b�w�=��w�=�Z���@E�v��+�K��`�;���r�M3O4�� /�ͣVj`ɞ�c�_c�,G�!W�u���+2,�#�O��d�m�a]�@d��v�������8�q�:j���������}���3�j�g`��퓻�7b,g�n�a~�~bA1:�6mA�j��A'��'�'6��ilՈ[U��'	�D􊲼.%˾����1�,���=�d��u6��R��!k#�۷n�cb.��nV�P����/b�EOf���+����(?��={׋xu��p �,ռM���~�N�7���c�_�D��r�������Yr�T}Op�~�6`A��kC4��� ����1?����c�U{P�0�u���"���}�ĸ�m�L�۰�4�&��]t3ޒ1�|�2���7��@A�lo����59���,}m#� j�d�Q<��^ʿ�A>l�3Qi��勽����P�}M��2��T�4o��m���O��skV+��/�Vo(f0��4���}��S�w{`je�~J�4��<Խ�E�4�rƾ�9&�GZ����T�	D�3�w6�{��1B�<]1p�N�������5�����]k�G-�`�O����NbhV��dlⓊ�!�
���7ܦ=r�9�Ki�|���Tޭ.��u�'�f���Lf��b,�ߘ����L�Z��e�ogE��s7�}�#��~�<�H��~��5�K�\��S�wO�wR��F�%�}�;|�ҭ�u���\)�49���l��`ә�-�J�eu��	A5Q��]Q�@.���4���g�9���˚U�Z �5��!D$O�3�ܬƴ\vzv�����3F�ʦ��0<�T*h�@��>	p�(|&��;��8�%��[�,�uwr�+U	�M��e99[�+�8�~K�jW�kk�ț��8m	l���+��lp�A�Nd��w&����TVx��߰Ŵ7؍�%
)�QQ�f�!��u�,A���p�ŊI�ɥ�/V�q�8� V����'Nj|��>��s��a� �7���}��ls���rH�Ħ�~�zV)�Щ�%��6���}ߔ�g0lF�;X�$�$)���	��^rT�P�9M�K!�����8o�OD /����챩¢[���߬�[9㚷�:�'�b���nwKA��j�t��x����Tv��1뱰�8^��A��v�؛KI���5E4!qNT��{�����<�����[�r���<��j���JMs)(�}�NlSCXT�2�"fYJ�V͐�K�m;a}
�d�IN��J�jŃ�7]�-�O3c�T6Uxh�+jK8Є.`?@I��<P���iϥWi�db��@Y\i���O�7
.�~�=�9i���)�MB�E��hL4�LmE*�ɣ�s.�Q�4%�n8�OɮYAXF��5����^���'��,?|m��	=
�U��������~p�Cb��-�[�Xe	8�kf玐dNyٖ���6��(olAP�v��]C�b�oV����ot_ 7u;����'Eb̟�
��8�h�TР���Z��y]���i��e�?�B�(}9 lԚ�*�''k��\1u
�WW�
}ִ(�킵*׸i��D�'Qv���/f'J��[,�}t]�L������O���i�F���ݳF@+�_ghVת�ޔ�?=���?Y��.i
j|c����%$x�H]}r=���^�7��wl�!���i�'��!$)�ȥ�ٟ6M���i�~M8�h��4��ڲv6>��w��s�LŬPA���8��p�Rt��i[޺�i��D]dC/9��]�	�sL�PC���R7�8p)�%�G�$�t��/�"q�ŽL�z�do=�/.�阚���t%>¾G�!��u�(_��g��yb�SY����2�ձe9�p�̍pu���l�T��>��Qq�\��-?����T�dyD��\��q �,q%��@�����K�9p�=��U�&�*�)�nm�s�+c}�>O.���!e����tr� �@�|��!��:|�%ա3��	r������7�����Y)Ԣ'!ecs���u �W��j�*�{�(cy�#���{��Q�i�8�Š^��F�3���@�"����d}�7����4M��K��~����
�	��u�L�}
x��X�d!Z��hZ	n^v���R��nX`�cH���X�pT�:�62���Q �M>��CתK�J2D��Rh_x�w���Bv�f���:�):N����XV}�Yo�3��س3�F\n�!nQ�`��C.Eas�G*��cu;���c�J���'9�mjt�0W��͑�趥�5q�NX��/���t-}�������P�;8�����N�%%���dtҫ���\=�On�GCX�/�3)>������A\��I^
�(���g��{��ֿ�Q�p����AJ���q����-*���3+�C��rY˖ �T�[�9����8�w�����4��Zbղ��榒����j���ڐ(��R����jV��if���;Ra�@�m�����0�;Yt߆o�^g������,~b�(�Q�0��~v�ӱc�D��[: �RH�́���	�`Ƥxo֒�w����t.�-(��$���~:q��M�h��.��bt=E��o��~b#Ϸ�xcv�.���L$U�dY֚���Ǳ�-��8����o��'멳 �n�5�ƞ?pi��zQc��H��f	�m�Eg䆄)��s��n8Z�+��#��o[�&�+fj� ��[���ֶ�4�Aq=$�1R��S��,u蔗���»�9,�CS��~Gs�q��Iْp��k�ׅ�e[o�8u�-�B��)��e��Z~�r*m��~�S�f�F�`��W�\�	�U�~H_�U!*�m����Dɪe�d��k���([S�9�����[@�o�G���;��Hg�N ȏEЭEK0^n��G�f�zR+�����a�����\�8R��r�w�o�A�����k:�j�<��{�;�i}Z]�o�m1d[볺� [s���g��<G����k���r�"�������[$��������~�Q+V�(���=����end�S����z�����,X�	2��b�
�����R��.�E)��
�M9�ӊT���2�&'ח,��`x ��P=�C�^Y�wk
�����@�pm���zf�8�Q�,�9X.`s�^\ ��V�Vz������:�8�]��I��`��L��K���:����0��o�s��଎4�64��۽o�:U��#Y~��w���L� �m�W-l��4��Y�>g���/	���г�^j�m��mک�eHHk����a�F���|��>�H�0xv�����%RD$���D�p]7�Ů9���%q�˒6��4���z0V�CU��NOc���o����>RF�My��a�܉'� ��'����{�.CZ���ԽE*?��{�}KaF�6�<}�7qKb@!���������-"�� ��&�jň�p�;e�����nR�ϧ6O�ZH<���y�8\�V�mJ��_��4�,5}��($S�gw:s���z5^ǫ�pGDy���0v���j3�{U��􁻆9��|<i&|�����Ρ�R�{���v��e��Q���g�N�3���S��h߁�(�{%��	+7Ձ��<�����y������G�)6m��R��.��4���I2p��U=��&L7P�43{��C��w
r@A��䀀ϲ�����W�*�Q���npDZ��ԉjA̓F~���u��43�u`S���|]}G���a:*MV���?�b.�2)�Lq��vY��HI���sBGH9ס���긱��jZ����h� ���xS(I4_*0�cmx�m]iߝ�A�79CrQ������<�}Nui�a�ef�B�L��yu�j&�v�gpoT7�'d\	6����B���Zkz���c}X��bR����C�o���:,�� �b�Ư�l��<)Rg�Q���z��@� �с(�?���&����p����w�4Ķ/�,*8�7�Þv[O;��3����|�� �2�\����`d��/1��Y��cY���$N��Ұ�+�-�)ױ9��k��%�쯍X�3�ħh�J��ѯ�#O��g���#��(r�*��M,���"�n������hB
�[�0����N��*J3e"�@�EY[l��4i<�X���l��S桧����m��q�$�"~j2���)M�V-hm{+�\>� C3�r'QNy���˽�o�%i��Uղ'�3��Ɛ��?">�
d!�ɣ�=�#���W�ĝM��Z�E>���sc��8������<�>->��i�H�����+B�Fp'B���b�Y�O��牲ҽ�3b����J��F�U"<��-�]�u��Z��q%����C���ͲG��柺�bR#�!�P�����S�h�p�
D��u�)E*��y �2E��YeٔP�R� ���c�m]��GM��u���nUy��	�rK����9 �FM�/��:��v�UwQá�^���/1p��*͖ ڍo���>��m�(�(���mF(
S�l�$�krWq�A�I\∕�������C����#��&���j�snmj��P,ɲ�P����u��j�Hdy]L^|�W�����6l��j6�ev��Q��JU]��2Jx�kVAP/c�Wi������	��x͕�~Lb��q�C�d���V�|����6e�KL(��u�5 �UC��zc>���	��\TX��B��b�r��zB
�H^��e1���w	{[�@��B�y�2���7�qw��9���>c��x�;D��1	�%�?��6�s{�+8��-X���a�(�N��g���!��򌻕��t�z:����ѝ<bG��J_U��q��?W$����o�����.\�ಚ�_�jǍ����>�����ޘU9�eM��G�! `���ZHl����3��l9�Ҿw�G�������'W��xV�wNZ�Rł�vyf.U2{�|Œ�U������`La9[�{޼�[���5ϏW���Nl�.��-�M�z�oo�9�}���#�ޤ���?r�^V�qk�K�� ����Uu�l$E\��z+ O�̘��}����
�����E�P���JpM�%�W�m�Ȧf��T��f0/&U�'gX�(�����Vj�h�_0|��jŕ���]\P��H@���x��|�U�L���p�$X�Ϟ;S��i>y��ð�m�/dڻN��Ff�I0���j���[�!O�?�d��aԭOlR`s% �T��T2cV_�qr�Ĕ<��óq��1_Wb>#wxt�׽�W�
>y����G�Xz<6�|��T��8��$RU"�*��3�P&�]�v;=�}f��d#�Lx�W��-n�&=�!���ǅ\E��	�ڼ�S��Eâ9[-ۉe�ZB��Cc�9ŨF��,E���l�<Mr��0 S&'v�yLU�>2w�Y�fX�������]��]���y�]U�D�!)a�C'j����
N :����ұl������(�͓^�Ӭ��:q����.��.����(6�QS�ϞϹ<y`s���H{6��^�K~�Yk�9*�қ5ɹ^N�Iߤ��h�
R&�~~��r!�)��c)��lǊ=��Bq�AI�9T��F���3]��0��f11pj�
��	�+z�ZN�d��8@=���_^���X��C�G�	v�d4����H�h�/����|��f�C3�\�m�JHX�8�m�d������I��y@e���<���^�b�3��m(F�Ux�����a�&�Tۆ 9���J2$֌�y;J8Ncv#�.����5~2>^�P���7r�cTl��uYY&�O9�����l6������@�~�h`|��qE�Oz�0��!C�?�@h�T��W�<���M�����	r�hv�֗�Ndk�mmjQ�ۃ�+1��֐��K]ؽ�@jb��c�?e��	\��=�(>5aK��!;����y�r���9��P\m|����6c�B��:�H��ޥ� u��	>s�<�9]&�j��5ܰE�K�g��jǲ��\|xl�_Rf����]p��gb�	�Da�8W�93���Yh=_����K���^�"ؓ_�I%>��w���V�a��<#+��Z�ξ�@���tbA�L+��x���H?�!���i�^�v!�C�a%�q�D��PQ���$���|IeQJ2γ�����`��;Q2uf���Y��^��w��3�1�	Qm��>Cңq�?���vyDZ�U%4_�'d	���p�<��������E���	����/�;���7Fb�H���6�a�y]�'�U\���X�vpc�������)�6�M�/[�U(�:���|-�nt���QM�_��fB��؀��t��w�W�sJ��o�)�S�i�z\V�|�)�Fo�1I��O ��L����4�)�)
���Ѵ��.������'���:�>g��b������n-&��7���_F-F~:����6)����x�}���p����uU���tv@"Ѧ��#$�aH;�a��;h���@��8�[���VȾ���1�u6�Nh&���U���*},��F��c&U�U�x�x�J����%���,vnr�<Q Y�D'��Ԯ�?�!�P�����ƻ����7���>�>?�'Lt��o8p;���u6j,^-�"��פ8�~ݢB꿵�az�@���/�,�h���ñ§��-�J�^Čw��}�C��{
C���>q�����x�e4p�UD��U�C#�Cȷ�emvi��S�\���i ��}]*'��t�n���-Ѳ�e	!v�
�(�n	X��I���:��Kad���\b:�:o�׃%������Q@6/�;uzΤ�O�j8�w_ޒx�*~9,Sq�9܃s���`�1������~��g�ū��o�&`t��C� I��6j5�L��P���h1�5I5�?S�L߾\N�^���*?�/󣯣G�
d�=9un���"��L�n��J֦�KP�X;�뾡�#ۍ[S��#eU�
y��T>�[�=ʪ%�=��0Ż����&�����R��5%MK�Ot� ��1�Y{2_e�yx���3�xl�7B��p֐M(��{�7T �\�C�ܪlA�e!�\��30�.'�.z�s���6�T�u���&���D��J|Xs)���z>����:���,6o]�fd����|�4�k<?�N�S�ƦY�<ˠL�d+6���,������J��Z� �}����'���|+R�dw��j�������l=��$hx6��V�~�{Hh��m�Uǈ͖u���xK8�GR�c�,�s8NUl�K�C5+��ri����[���-x(��u��,&�ߺ\6#�	��@�K�jy��h!�~�*�2��:��Z��Y5���j$D0�St �_�D�ΔR�x���� vT)q�cOG�ܤ�r��%I�!,����U!P�/�� �8��X,s&^�؃�3�?)��0x[gխ�� �\L��R�F��Z��W.�v(�r���:oߴJ�F*,:��26f���.mX�Fb�s-��f� wol���39��5�)?�"�	�4�hh�Imf�>���ZV8ht�-&W��?	����@Dz�������`�[U��Poi*Ŷ�},�Չ^�8��u+C�b )�!�BN�`��n�V_��o`���tM�u�	ڋs����|��:�̜�~�� �B�5=�l�}KpZ�r�؄ ���ib-ziD:S�%���^B���IB�v�f�P/��Mi��b	��>�U�C��.��1:@�E!�Ijsp�L�)����[���`+�t�`����.���npI����!yα&�r7ˋ�v9,���5��Z�p����������Kv�ٟ��RZ���0�=�J��q��隬�"�2E��.���/�:��]s�y�4zS�����~��-.ػ��?Y��E�[%���Ma2���~ac2�����d#b)�wӚCה���2`43o��R�7V�sĆ|lQ��H�w Ld�(��������b���䴂�弙(ֲ��U}����a���&��L3 ��!gE�<�J�q(��V�q�}�`��e��=�<p����o����W��,����b�- a2|���rk9����qY@�@\r2�r�4�`j��,wR�8����ny�/9�J?�c��9 �=*8�Ƌo[�p���T��7�QjFH�6�չiaJ��N6t����֩#8��oت֒H��`wUE����Rtp�4P�y�:�8]���m�~|Q�v;��X���c���Hc��x��zZ��ۚ,����a�, �Ә�TEe������49>������M�U2�7֟1��B�}�v��+NA魝$�bD#�Ck�NG��$��@l�k#E'v��ˬ�$��4��wh��"��2����,AC8�͑S~�dgꏮ"b�5��U.W�z�I�bת�$�s6���+*&�Y��q���*�(2"�ˇ��f�6�ކ��쏗�*�+�RG#��{�������a��D��~3�S�S|S����z	2�$)�����d�E?�J�[�q����
��ٗ����Н;	I?���w���.���7����e������C� j�>��㔸��n�n$�=�hqs6�S�`r�N0*
�J�١"���A�T(VG��p�i{g?�6)�-/�ڬ\�hGh����7��k�֚+j�����)=TUs�g@�J���:B4�t{5e!�<^���gԉցsz]siN1
8<�s�HW�~����x��9Z���<J��bz��fd����b!��w�
g{�p�~��a�R�����~���jRp��
�`j����:�}	p����}�MP �F�M����T�6��6�����|\�ZuQ@�ͺr8�/!�&<�c�t�4)�����Jv*�5����F�	��njc/)��W��@^#�'&XXQi[xy��)?�ѫV�r3xG���`�%�����)��xВp�����;/(Α6X~O6�{�9b+�i;�h���b�� �d@�z�p�������F�G޴�s|�/�E��xr�j��Q�'�Č!K��\n�!��ieq������Q-��v�$eB𨍐����+�d�M��
D��]���})��V[ �Q������B̵5V>%I�zT�o�ѐzӅX�Q�&��=����,԰����@	_����F_�՜�n��o~!��w��y���\ГS�8e;:��T�T:�h��W��9(�H��M����J��>�=���Y���>0^�}��6�p?���и���H��x��.$*�� nlA�q��g���,�'�	�ӻ7P�w���#a��)>+xB��x��BT���Q�L��l���;�L�w���߅�n��פ.��*��������,�~��A5*����l�J�F�v�:Լf�A�$�9;1�|h7!:�j6Y���NjW�Q�B��u�w��[& 6� s� �A)g5Qy~Y!e�Pח9{�;�qĦ��@I�[��v�<�ؿq,>�`�v��6������u1����#�s��{ԡG<���^]��,����xsP�w�t�s������\�tps�9�m�i��[~�h�=�򍫛��rTA�1�*Ϛ�{Ñ"����`.,'�KՑ��ZD��F.A�Wn�{���s�n�@bgЁ���Brub���y�x��*tp�Mi`6���Ɋ���,��ow�5� ��4_J�nɕx�Mh���߯���a/A���,��*�Ǜe�|��x��~�ī�!��a���$�?�l�պ�����=^e'�*���rS:�6c��gq��I�$΅=�` ��T�k���H: /TH~_T��]u���Ax��_ޏH*?���ǦYD���T�]e��<gQ.mtD�z�>���JL0T�H�6�XC�?o�H�.$L���B�U1��MiQx]��iu���4���纓��(fF��ѷq[����O4ϓW���Mj=_�S"������f�zX*h�HU���0�'5VP����#�)'6L�.��\��l\M�������l��ã2x�qs���1V�u�����`��j`���ߗ����:>MD�fYh�Y|�
^���Q́�[�I��/��b��k�J*���'��Gyn~^	��r4~5��*���G�0 E!pf� g��ǁ�n����y�
�������
�]@M-)j��+���i�O�e�����X���7n� ZtU��O��7tEWA����x���8�������F�\�j��b�9�%,�)�F���]t��5��I�Ky ����:�S�Vߍ�W|_�	�<�&��������˕��Xډ����ɋ��
CU/\`�ec�~(����:.Jw�T�LN�W������Ũ5N��O}f��F��[�c�Cx����.��I��NM�}��ʧ�y��_��qf�A��^z؞8�`������$�:�\�h/gx���M�^������E,x�#�����ˤ��nD0�b�����z$��׸�`S�S� ��N4�7(ȴ�z��������B@r�7��Q���V�ɻg3M��OPm�\ԡ������zn�������?��Vɧ�w��aH�fe�i`2䉧1
��N7�N�5T�kf~^�����F?�N�*.G`��v��cdq"�Ϩ�&i5�M,6�񾶟�%4І'}���;���q��d�;�į����o����^:�|//���a��y�1�]?*Y����E�I�&��@xdmy��a~�ve�ϛ�%���CE<&�p��H��x��>���,jH�춒��c�r�-v�a�遠
���c�7����t�K�(l��k�*�z�+�ę���u�B�y�ABdaR����T;��\�l��(_�7�
�xƉ����%[�7�{@bs2��m�	��J��*�)��XB
����-�����E�&��<�%��oT��;��z2�q�3�����^�&��+:�#����pb9P6��w�E���,!����O��b���㼶W��(Hd�9���Zh�%M2)Ȟ��~�Õ�w�:�a���+�e$��)���������|D��^�k��U���M� ۽^���Ts�Je���J!��$vs>{L�A>��Hl� ��6�1�3��n���z����Ye���+�
��_�9�Q&��3�׹�?5O��n�ݭ��$��e0c[jP틁��*|�Gup��O�;�l@�x�f����Ѷ�y<f?5=�<q؀��Cw��k ,@Uh^pm��������I ��/��z�jf�#��+}M��ڂ������.�H�>�Պ��m��E���Y9�g�.ɑ��p6�ۘW�����[�^rif��П�7�Z�g�;x���WX9�$A���&w!�9-���u�оs���TF���W^ C��-�ڜ���Ż ��zW�U����Rw�?r֙������P3]�|��p�W�Oޙ�ƌ��n��~-~�HIxɅ�+#|]KHh�`�~J<�/�����
���]�k�:�眕}q[�H��ĭ"#J�D~�5�>��y����I�@5Rx��GV6�)W8�H8OB'� �o��L�(h��g)�����\RB��7��ۼ'2l��l���pf�\V�^�E;�~s����K�b���8���Z�bat�;x:���N�82�cZ�[W-�sˌ���P�i���1;	"��b]֎-m���idpb��bʧY9��������-}+ђҊ�ߢ\E�F. l���,�T���nxn���A>G
��] v�&�7��}�}�S�$��PXͶzꕦ��o"7��x[O>)T����eo��2�aP�H�ppH�P���bfvx�)&�j�Vע/2s�s ��MG�� �F��9�Zm�4k��
�ojq[��	�H��C��6#�/��k̠㇨E����v�ߊ���ߥ�����s/�p������E��j����lx�tQ4���)���s�:�!i�qC�N�v��V�Y�9���`�A��-�
ا�
s��+�q�ʮ�n�ub48��6-�]nP{��$�G2�_Q9>���h� Aϔu�8y���FD�Yps4S4:��_��G^�s璧�`����EzT��pZ�q�21���t�#�tf(0����6�y�}�|�<G'T"_�މ���x��>�C�¼\v�PA��*#}���=�:'F��䵳n�=Q�X��%�,޴���ĵDV��U�9}R�B��k�z�U�w3�|}�(3��T�!H6*[VԘ�O�ݻՀ)���~�7�����s� f$��O?��H����Ԇ��|^^�gf��3N1'/���]�T����	moZ�*J=�`���p�X\�Y��H�"�L��t���;�c���.��>��70]�_�����9�3�u�1�bW�rEcz�F*�V	Y:y���)Ie����c��:6��hݲI�����U2�#W�0�Wp8S��W�
�]���8r('�o�S@�hܣw=�����Gs��q�2��}��:_�Q�j2+Sk� ���:w��g�����Z8��r����>�Y]	���s O��h�$`�+�s�e���@�|K8,yc]�쵂�\@���P�`	��Xl|�)�W{q#�+�o�����Q�òr�^�=w�����m z�ߪXnY�`�ۿ4_p�"Lo/5,.��@�I7��}�?~ik�+�%]�N�׉l�Y4�!}��Y���aa��! ��4/���l����?�Ԧ�{o�]��D���4��*�?kSӻ�̺L����E�����v�m����Y��Q H��a�����=�G1\^�P��@�뱶(�J%��G"!�9:��� Jҩ�WLEc������B箤Њ��vj��0��
���k�A��R�^T��,����"U�n�
@�)N��m�K��UJc�+��G��f�Q������-O���s�O�����rۉ��a���I,�����Oщ�e(9R_�*�g=3�x�E�6���Es~ �p99��IeX!�btM�!�U;*8��U�}�,��ME��-�/�3�y��)
�f^�����#� kg�V�@t3���A8�8��h��-\?\X�/�D��>���$��(Ұx�.5�y6�8|4_�w����f�����#�<�&�'��ۘ=�m�M�LY���r&����l�����S����{Be�&�]^��e�P(v>�"�e���Z�'d|kӈ�푐bN'.kA ;�ASA{�e���Ú)�Bޙ9[%&����Q���Qȓ�EU��#�P�e]�D�[jJe�sJ��Kd��f��3]��Z��RdG��[������p�D�����x~	3g5#Ư��j���R�T� �c��XOĤ���X��9� <9v������$���ǹ������O�N�E��mح�N��������VL���jH^��}1�q Ye͙>�uO O���>e1Ӎ[�h�[n;�i|�}'�٩���B�T���UJ5}lV�́&���H`��Q������p���/�00��!�)�"k�a#F�*W]r§yF��(�º��"Q�rL���0Y砰'�2�/Qt�ź0�SZor�A}l2��w������7��8��S+3=,l��@Q"_l;=�]����C��^N�Zލ�
�*8]�X ��٠�y�9M��8%�@aFd���F������=oԓt��̘�B�*YgF���V�$2<���)��;Q:��+6�N�
�V9D��Z8�J��W��Mͬ���V�b�߮t��~�vG�!Q�?�M�f�b�a�~��Ku�ꊩq�L^�ݺy�j�>��1���j���Ҍ<�t���e5��sz�e�j�+��GP�dc��m�Q�_:��T�XJ�,�2�K�֓��o<��˱ԌÀ�_�EƵ=�/��o}Z���kU� 8��#��b��9_����]h�F�tq���WY>��'L��(��.a�ϠʣD�*��ڨ��|j�ୌ�UV_]E���^WqJ�x��3`d��b)4$rML�~F_�:mGT���;.T;��>a��f���1�!�M-��ou��P��9��#��6���0|�F���$Br��s���ht*KG�D�v�� %�=��/�՜�k�-���]R�Q{܍Y�f�;1��Sw�9St�/if�=��6b�0�����媟�]A6��y���,���gi�����z�39Dt�)�|���C,<��>���?E�:�{Ȍ��hYR�]NF���4�C(��w'�ژ'�c�$舘��oi��m����o"�-��[�!����j�և�J��cME�N�[N�lx: ^w;��=c��93���`���o	A;\�8R~�`uVT�ZkG��v�w}��L�<R���A�A��H�qЋ��f"^�oh©�j=�,5*���\��v蔬%H �a��K�v6��PI�[�%�+��[ԙH
�������gy��U��hH ���6��<�$Ŵ�#BܗXD�Y�L��i$��FSP�Rqd��	�.��z��q�K�n��
�]giJ	z��/p�v-	L�a\|��\�@@���ao�&���c=��2Ng��i��`;����<ם]L�58MP�� �aC�eMdX@�� l�E �`��Ȯ^t��d�^��a%�B�F�;�z�|m���y��x4Q)�~-�*Sc��Zf�oe)���
Y�>6?�:_��/�ˍ����핛f���ҝa�Mi���J�\���&��WAcup�#�`���[}07�S�	�d��0����@v��O�]z�=�/�+vQ��'c�t���3���7�ZϤz�m?�{yϒ��@�oo�k���M�%;-�
��� O:������7{'�7o��	��;2�F�h�U�|q��j3.�m��zYs�fj�?��0qM���Jy��z��e�\h��8�ׅo����P^ۛ��&�?u�.ʳ� ~�d'��o͍�r�w'N��?�l�����0��#�o�.�3$f��fRH|:�R3��6��v����r���*r��c����My�LMwf��D�X@¿���]SAS�$O�
�L�Lq�#zz��Q�	vul��A�-�6C��A^��.�%'�qB�5�e/��l�-�L�nQH��ѽN����۵ +���� ��S�êL�b$|g<�$Z�Ζ;�O�����)�pN0�ϥ�A��P��g��^�Y�/�}�%^��I�bm)��^~�60e���U�[ ���S6�Pk�W�H�Uq{�����bFBG#�z^oL�~��T�����2ݴ���Y4 
B�ƈ�L��]͙i(s��pT9ḀcL�t<J���#c9@���N��)Q� �ѷF	��|�l�[�C/��KՐG�D{m(�c��Q�����#��{�D���
�1U�VYAkmfD�@����������G���M�M����%yEf15[TQ�`U��:,"��{,�0�����R�[�%������J0�� ]-��h�ӂ,����3q���'�Vnv��ӤN�o��Rb�./Zo��/�R��.��{�i-A���b�\�t��<ǌx��0�ӑ���.¿��^��w��GL��8Q�Tq9N)*qW��I�g�I�c�r�6�����S�\�c$v�
3H��q>3��d/L�U-ţ�!��qq�F ��5%�;sh���z���r���D��Zu��o��]���a6�*ZrHq�J/28 <S�3�|
�dy��~f6K됗>ږW"mpm�B���,P�[�������'���m��\��*}�OO;�Ra���޹8�0�,rbi���B�2x0@J���Ŗ�c��(�ES��4�{ꟖA��][����������
pF��Zv�b��*>��Q�G|n�~Z�@V����'� ��H&D/�)���~Q=�̗n٨Ͱ�{��_Ҥ�a��"����$�R@:����mfEs��=�}8��5?�6ۢ���8�C�o���X�s�o����C^J����]�oZ��p�ۼ�̈��j�IY��þo:�����r��
M���m��6�%��n�O�g3
_�Jǁ`�7�����!�	/��j`�����M7<���	l�@�#ə��	LX"����S����'�L#̡"޴�}$2K�	�:��L ��gkVPbut.�|���z�_g�@��҄f)������_�Mk�\�R�)
�4���K!�y���"V�� ʬr�:m+X��?KڝT�-��h28��d-��ۊ�d�P���eL )������cU��U!�v���s���h���o�����O��VFZ����{�Y<f3 ���ni	z�F���H'��7�cg0��d��Vw!:� �v��!���2�� ����s��Ъ��?I���4I>����pT��h���2%=F�E������	T}��}�Jҽ��`Kzؽjk9�;A�b�?[L;�S�9<�Q�6�<c1�3�~W�Bk��
�'k�;[FݫR�n�y~#s��0hh�P��5#�xG1Ŭ��ڻε�ȹ�����ue�f�% ��G0ep����ˎrr��ó��e�`��Pv�� ���X���u�9c�?�ٜ6����}_t�%Tv�H��Ex�V���-�����:�b�ץ����ə	$���q�rN�fPC���S$��]�)�|d$-R
��聡��T,u���8����eZ� z"�u��u��p���3�����K��FB��X�X
�n3��R��gI�;�5����C�J<�ܧ1x�;�X�QՙY�W���N��D���P�:�x��#c-������&��2�vo��tSxn�߾��(�K�̰�-���&���� T>jQ�fٰ($�;��OBR=��I���c���!`���?s�%�jP��R����Wǒ�Wꃼ�c`Zԗ2^J�׉�z:cYdsq�<�b-�!(�¼0t���8������~l�}~�E��[{[�q��U��T�Zc�0�;�
�~V�B�\�G�|�:��=����/�qix<}{�OlA]��pr��<��/��̠[h6 w�D�"��va�����Ǡ;�=�I�?�J�;0]G�+�`�����1�<a����La��ȏ�����ԧ+0�懶���_����1H��Q`!iX�ʇ���*�ί@Z��&�w��n1mr"�憗)h���X(t��0��`Q���D*�
ˉ�M���Y]���i��<M:rX���4�R:��N=~f'IC��|p;4t$P �о��Zr�U��i�V��M}���#�����	�D�b,�B�Y�s�9��_?�����F7��=1;N��7o%�8��M7�L���]j����_��/x�Q���}�o{_*�t&$���ؔ�r$���?��E �;��HW,O	��|�$�A�,-6xor{�j+�S��Y*���� ����j);�7"t�(����6���G ��g�K�M)N���\��Q��c6ap���a�5��+�$���� n����J�j��g �Rh�PC�\JTm��"V��i4�Ͻ��%�>q��t2y������3�Dr]��|��[.���|�����~�o���~�̧�vR砏Y�h��dNZ�Q6V	�iZE³ߨ����4wB���:�g`��^�]2*Y����:	������ܮ��D��H�ZC��P��5�Ҫ�GF��d��K c���9����7����rr&ea~�nw[rty��eGGK�-�p�o�n��v�?��<��.����!���!�$p�r��9�D4�X��fSR�Ml�����yO�͠`q�ی�^�k/�5�䣇X�O�/D�'6}K��>;�3[��h�@`�2`�J�P�HK��p��/��-��)��	ֹ�ꑯ_f�u2���כ�k��W}p��|�D��Ֆ#8��je��B�T��`<�Y�؏���>�Fh�F��o��v�{Ԝ��%��д�yr�S������|-�.���2RzX�[|E�D�W��܆@��,�� n�E�u��8�o������x�GJ"u����uO�50s�͡^���c�6�{n��a�o�>qw�~^)A���xoo�%V��7��"�]^���*��CO��6�nԋ�v@��L���,! a�z��ڨ8-g�83�S���l�s�T#<�E�?Z�^�������b�A�hx��������q��NbnH�A&��_t����Yjsǈ��7.�z�t�Ѹ�a	�ҍP�Q�s�ZhK�M ��^�[��\�n���4t>��I�W��xɶ�O?�`<�?���7���r���0o�؞���Z(�դ��j<$�c��@G��&Q0Z��B�Df`Y��M;Dr,�X�p�<)�a�	����銒�i��6%���ּ;�U�6�^��"�'����E����Ɨ��4�z�<*�Ӳ���o��dN�����Ź�QG �A�=��Y�����8��+��2��7�퉮]W��8��Hɜ���ֈ�	w�`���z>��{z��F����S��{�[Ԥv ۉ7
_�
H�zȅ���p�Fl�!�����؋/��e:��m�����������A�5_�n'}o4Y8�����A��1Q�th|7J\*�ڒ{��W��}M���N@jZw�x��j�o��"���7�� X�|�A{�K.?���G������oU��h�Ph"�לp�k�2}S����^I~^x��ޭ����2|c��O���3é�ڷ5r�4��.̀��z�S�����l���/�ZkM��!�V���%�2�L|իl!����Ե
 �h��7&�nv��N�#���ǯ~�u@���]�QEo��?�ʂDXr�Wb����� �q�?�f_�v���H-�끜m�4<y2UN�-h�[�{���!�F��gn��^����yu�`���}����[CN����Foa�,3�[�f�a��y�΍��<%�w���K�ރ9�%���|B<KR2����m�?s�2�3�XA]s;��p\0��g�J�C��JMAv�v��6`s�}K�՗d�>ܵ{F�e\�eW�^�{��є]$@[M�V(ۀh�����߭U���I~�<z)�F��4�	���0��ܑS��׮Oy�+�]Fln��
�+N�i_�V�0p�5���XO�E~�Dw�f�SvP��1R"*x��0sÌzW�p�M��L�5��|�!t��C�"k�9B���g�BцX�x��
x6S|ߑ��g�~O,6��
Go U(R�|,�@[��g��� �R�C`?���2rT��R�u�	�ONf�Z�0�IZq@9� �U�dE}]�u�>:��2�Q��ы�c�*��<S�H�Z�N؎K*�8H�e�ݭ��/��҂�;F���٣���7���!��S��uz<Iiۗ��0��1�
��$�Yyb����lw���D� BTc�?(�ry�"�V�K�{�-�?�/a?�>e9�����f�fX�9 ov�_���T1����u�ײ\�B���ސa`�����1���t֮U��s Ɛ�#�WYl�'�ĽKc/S�&}��oٺ�w��� �����ř�!	�4�o�ؤ����/�y&E/^#��Fpho���GC��Os�2�{aG�W�w��0�~f�H8A�+
v�����<xw�ºQ4��M��b���+ �B�V�w.��C�Ԫ�/0��!l��ꠘԷX��ƘH�
�����y���m� �}�t�c�+:�|�
r���n�v=0s.IL.i���:^;��-M�oKCZJǾ�hn����K*�¸^_P{��5h�SA��I�Y�0�,vP�;���u@�<M� ��,���Ɓ7�w���XǮi���� �Jlŵ�-� �ʽ�U懗6�X�x%��R����9�H,��A-Bt���m�螣�X�3�h_>���� ��lB3G�OK؍��3�\g�������'�,�2�jLIr4�q�j$���������)Ұ�?I�RT(���d%0���}�4�Ww$w2��UO}�B@�򄨅�_D�5�x@��E?E�(O����b�����YG�D���"�M��<���!�H	#)K����܅��,�,�k���=�\'#��wR�
��[c�"�4qڃ���,�f�޿�%��^]e�L�904�ҏ��'����|(R�F#�Ǎ:�}	�����o�f��e|���m��d�L),j�8���ɦ9�D�M5'H&v�S:��ϸ��A��yPUbe+r!��J�]$�ֲ	��v�ȏw'P�- �y��c�O �c�)�����vj��!t�����������Q��
�Ӑ$�D�p�%����=�d��;�k��*7�?��/�*�
Nlh~�@�j<sQ&J�͘	�sѹ�ց|!=s���5��4�.� ـ���d�d�P3�hڬ\�����N�no~���j��\dq*�d_��V Z���~��x%�f0��`ķ�v�N�R����Psg�B6q.[��ռ���F8,H-4�nH��-��2#�x��VB�*��ݦ4��o\SR���{%F�aK�U�>A�l�Z�q��1
�<�θ_���Ѿ.!HO����T��Or�Bfx�;$x��錠 /�M���C�R�s-~kݜ��@���Z������0��%G��Y?���t[:Fhvh�NF:O�̴��K
h��k���A����ӱ@�YH��!�A�BO.}܇�t޾�b����*c�˒RA/�@��7�įd�ԭ�g�dT�r�B�
�C>&~�ZN�*�]Xr�ZtG�I�7�'׾��Վ�TJ�MS�讃�����5u���v0r�?T{��?�u}��u�d��ʯP��#����q��?�Sb�H/��O������G z�1�e�-���	���e!O+�#�ʸ65�ޱ�xu�N5�s�Xu��U���@d��aH/�Ȃ�t��_�;�"R�:n:����?uYN��]%Pw��C���հ˗��j���A�?	�Ǒ<�M�!e���8�X��|��.��{5&:S�u_�R�Y^��hֶ���gz�Z�w�0F�':g%��~o>�Ld�L	�׋��{��3p�/�₮���G�=eM8F?nueI/ǙPh�s)w�l�|�N/v�A�V�P荱��7��o:����V::��%j��}�!{�����9�i�O#R����J�;!�����7��<��Ӵ�m��:<�KU��u�~3����^�!���|ʋ `&�'�flA�� ֒]C#�n>�p?�������H��������x�IJ��X�(L�fv�WZ���I�paW�Ța_^�f�is�����0������_����Z�������Q.`���JB��K�s�Ara�(1n��[��y�9��Z�<c��B΃:Y��~�M���t���+0�_m��N���� �l�<���X����Α��- $^-�7��9��TRQ�@�[�
����/��|?q۟��֥�m��h�"��@nh�>��)}% Ђ�	+����0a�6yd4�9���Pf}�Y.�ğ��6:`�|?6����c�u(��<w�o屻����;�r�-d�a�q��Aa�{JmJ-�5K_<>�bc\k�R5`&d��X<�R���.}xE���A�e�Ԛ �m
8Dë�d���n_W��F&��恏Y�;�"V]
p�6于��#���+�d3���D�t���z�1�KK��yl���49 ��8f���xnpr�)�å������*�$B���C�|�ƅ'a�y,��G�����يC��������x����g�ql��:Vϴʭ��Z��q���Ȇ�mN>��.*}�:��/ �I��l�tj:Z�A����ZBøM���k��f����9�:dP�e�۵���-+�RU&��Mͷ�r���A*v������Q���c�y�(Ʃ��w�5��v�/}�p�3^��zMuK?d�^rv�]&��b�F����'mB4[;2����VM�	] %��;5c���Nx#���Q�?밵����=]�xCW��䬟�^�(�W��o�Jz<8��C��cZ���O3��I�^I("��"�=��v%Rز�����I%��j7%�>�HC"���W� �H�C�z|���vG¨�:KK	��Wd{�2k#>��7ʆm�J\��ɲ��6rI[�:׃�I�H��T庝|.9�����Ĩ�g������.!��>D������F,��p(�G�a���A�	1��s�(��D�{��j���h�u�*��G� }@���k�|A���� �;�'_O�+���������E&�G����˯$YY	$!�ꧤ}�C����$&l`I�u��R�FXѮ筞�r0  ���n����7t�X��~\ʙ�:Hf�:��4l�%U�q��Q���1�Fɦ
��&��@�ۿh�����U���OR�j�ȂU��4Tmیs�ţ̅,utM����.N��)��Wk���c�Y�vE
��M|z?��`���b�J�(�Q.�([|Rb���v�b�q�E���p�F�wZ�?�^���½H8��/ޫz8I�l��S��o
���S��g��ulB��	���CYn1yO�󫏐�d�_�p���ˎ���XßN w�6�1�z�}�+����+�w��ri�Ą����B��HA��a��	g�'{-��7�I3Ƈ���\WG���o��c]���oVxk����ρ����� �H��)��=I~�4��qE�w	Dv��Ǩ5��0�Iz�E�?sh���s#��vV�bﵠ��N�ן��[z?�Z�z�ގ���=`�ڣ ��Cl)����W-}2UWs��ʅ?�QC=-�� E[!=TI�ϮI�q�MB��aj:ފ�5P�`�U����b���~R]����l�R|��<"�z��|�3�9�v\~�j������j��6@ry����!GO\�c���-�׆��i)t�\̚\��_�<l��WK����(��'̿�f{>� r)T�c�l�k.��?͓�n��&�E���Z���X�~��s�����A�3�	9,a�[^��-�)�I�ÅI�Fw	�L�(Y���46o��`��/P���]ȱ�j=3p�G��Mҙ7�v�T��-Q��s>��>�>J�<��~G�V�e��G��u��� Q�y�rZ<Ј`=����Yg��k�B��<,��ʬ@����)���7��q-št�Z�*Zѧf�6Q{���c���� ��R���|�b��;�.�'͗P�R?p�}8� ��l��|4>��q���e�c}�,8��83���c���]�L��(�ɸ֠bw��9ף~)>C(F?�@��t&[^���$0с*��7[*P�=�3�̖	���������@B�E���~V��K��L!���M��6+��(/g�KY�xj�J�ƣ���7�k��%�KxIi�E�ٿ`��ac9����th���
��حs������m�K!	\��H�f��}��Z�@$��c�'//��0M�_���G��Z�\t�h��gJD�e�ީ�3��l�̕gLi�c��lAպ=H�1F4�l�H��[1��H �؃ml쐃�����%�u��L�N�[��P�����4��e���e�ǿ���gc��S��z]q�f��U~O��m.�=�_���Ճ���g�N�2��f�.��l�hQ%1����^ӱO���C�1oL����O;���Z��Eޢ���\0�u$2�P������y��R���^�"�b]�}�6�3���C�J[qSZ6��$d�!���W�d�]���j��y�*#�.#V���F��x;i�W��"�2������NH�-���E�K��_Z������˳�����9���~j?���I7�uM�yS��G^�ͧk�-$�L�.$����2i	��g��sFmM����%Iʔ~�"�t�����ZB����8�]�,��`��NΣK���y��j����ܼՊ�X���c�u«��*\��y�uZ���mu���u`>FB����Ji�Ͼ���ƅg8�\�0H��������\�;	~M���%��@����v�Z�"
���
" ��}q�+U���I�M�'Ϯ�e�v��U���,�'W��Y�>0�J0�ɡ�5<�8�6�ԁ��N�I����\$�QI_���5��������e��iv���Ť���e�ܯ�`M�M���)���,�7ʰ�	���^}kR5�L����%[ ��O�P�Q��~�����JS���7������*�� ��� �+�h��i�]/L��T����̷���O84q?�byh�g=��ͩ�25��e���#U�_DG��#B�/�o�:��{-���)�������5��8X�����I�o�ͪ`�9J=���|xWƘ�0 /�q�%��2�W�7Hz��ΏP~)'�i<�ڬ'�id�I�Թ�2A;���y�-�䴠�I�~Q��?cD��I��"0�0��F�;�����v��o���CS�ԯ���l��|a�û�?�Z�I�����e6M���S�xܿ�����q���{S�C<��.=_;*����:rXp<\��f�h�L
*��2����kD�ԟl�2ݏl����H�hw�wK`�	l�������|�,�*�]�	��F���!��8�B��J�!05�I�anN�3�6(@ST��/��"�y�L蟔�m  ���ڒ�Iuг�m� ็I����̓8v�ɰpQ�y�����?k�X�čq��~o��#�Sx�!�^)a)��BI��>�-p�1��ܝ�%huJL�d^�߱sU/y��hUgM���Qj������Q�(�x��OЏ��v�Wz��GUDҫ��*����5�h�'�u����][�G<�"BH#e��
��n�ʨ�����S��M6n�
/<n�{��`�m���pP�#6镄�g��05(G���̾��-ox[��2��p�^$�x�<�N���B�+�5[öfĬ��2��qWML�[
rЉܛ�����tb 7����\q� ��34r9�+���gg���@bS��`2JB-š����R5���w�.�C��Yu�P�/I0V��K#�m~T3S�g��c�$g(��h_��a�&oF�V���>� �����&�I��zN��l���|��F{�Ar���L0U���?����p����D�_�_[���U���(�J�G��(�jxޡn��(oP��Ң�,�wԇ�k��7�@�A��A��y	�U����H�\���'|���/��k�y�*��Ԭ�*T�|�V�
`Z7)��}) �/q/Y�ǁ0�'EJw�j5�~Y(���D�7B`���ZJ�

��w������>TZ3�L`!�iKڙ�+Mұ]e��C��\�\U��tRK�$�7��)m1����{ #�*��	?K�ǲ��s��e''P��u����W1ֿ�tGy�5W �>��J�����>T2���X��{)~��ui*u.�Q"�))n�H�jm����(ˎR3ϙ�l�v uUk>�w��-?\����;4��J��%���g�n5����N��dn��"u��Yy�j��z\�e~��MGuwR��d#��,��p@�J̤�P���Gt��t)�Д�L4W���s;������(�/i����� n�{��2��m�rFC�'��w�qzLGbר�@t(Z���L�>�k^R���_k��? ���e��� 
�|�͌�w�=MQK�;\�����{f����~�Z3�.嚣R�c?�b"E�H�8u.�F���)X����"-���˘��.7[}�����D8H��Bm�����P�^d����aۤ}	cig6BQ�_9o-�Rk,9{
�D~łہ��
��-��E0B:�á��JS��\���1����x,�p����</���E�6G�xs��e2��^P�B)��P��$+	�Af@y��@?_��z�.}���1��9Q4K�ц��L����D���X�.�%��#Q��TQ�hĢTu�]��#7�(+Õ�B�c7����d@�(�jD�3�����E؉�r�ٌ2�w�G�(���*"+����2��$e��
<v�\G`t�$ޡ<���}�����?+OF�w�uNTG@��H����T`�K	�B"X�K�fFR9M�P����k��Q����4��o�f~+�������O�/FXy����VNv��)pm߬.'&x�ް�Aܑ�P6���5�b[�/�!�r�5M?�8"�HMm't�"��av����;�6;}wb�#�9k+�>�W�!�!� cE�|�>�B���nB��,,���u�D<�c1�YX�	D ��SAq�o�Ejpv2��)K'�����v��D0eg��ޫf|�G=2&u�~HB�v�æ�_�o{3��oBmk�&���j�����
��7���8��z�������Y��y�6���2������4�`;�V]�!�v&�b(47���Kڳ1WY: �ca6�$��k�d���&�e��
	�3�/�=�ʛ�	C��I�5��Ƭe�@�G|�~>��u�EӒI	X!w�I�/�s8�Ⱥ����v׃!P�k�'&V|+����X��3~0Fĺ����v$�~\&��46+~ߙݚ����T�S`�_���kL�!�T����C�L�(2�e?]o}�)4ak R� �.NpO���L���9�ײ8-3S'�S�;H�o#��b���~���-hW=M����+6}�ed^Y~��6��h�u������Y��^�gv�g�N��ZTY�Q�6�n����va3�º�L��hC�	r��я���n$�t|O��8����6 Ei�pyp�c�y�P��&K��o�`1��}�^���ģ����Q��a�m3׫tXE��=|x�
�t���.8������9��Ʃ�(�zB��|��^>�z�0�g�^�{�ˌ[V�9�l���� II߭c�sjq�������- �ʞRW�����#B��Z�D*0 p-�z�ԏ��ě�DG�{�E����N��­h�m?1��V���QA�&Y2|����Vh;<�Q�'�S���ג|"��<jnf;J���*�9ٯ,I��t/gWC�1j/ry��&Kr"0h(2Q������Ɉ��k~HK~6N�.0�C��]�2.��-7԰��J�lb���P�7�66�e��78{eJ�d�ʮ4��O7�W֛ �߶,i�t�!9i��,�$�;��;~n�3��t���9������?lID��5.�e0��sv��*.�4�V>��,�� :��3鱲/�w�p��׍��ׅ�'x��kv�U��(��)��C	{�{&E��5$By�z�v�b�ؘ����n���% ؊���h��S^ z�r,+����ʼ*?[��uK��T�h�KGD����G��)����d��}���b�/��.�&yE���s�a$xxED����˓y��m�ZZ*G2��Eޯ[�%����)�p�>%{�L�����_G���{<�liKt��&����Uj�B��ҧ�H������3[nY�ledh�l��:���3�����o���b� J.�DC��}܇0	�~� ����F*V�̯\O&����=�:�����1�2g4't?y�$��}�m�~wI��J�����S6�k�V8��f�CL�T��P�xGh�����m�Y�7����~�������随5O{n���ν�g�q�K�¤%�`
O�� rR<���m��Yo�ڧ({�Ѩ����=<�
�\�����tv���3��
��n�]S>��l����{���p鹍!��qJVҭm�_]����B3���B0��:οo�۞gs"��.cMN�4�T�4i����WΧ(�LejBS�{�"�Z(� �|��SVQ��9g�KiIk���P6#O��� =�9��|��Q��R���x���Kt�\��n��a�|E|�vRe��]s�gK��#�B~@p3噰$�ūBq����M	[�R�H�{���TֵQ��$��ڵ��N =k\�!X3FZz̮��i�~c���Y�d��W����/�c��1��mR�d\��Ft��ɼ���@Q=��������Xc6%����c�B�,�E�����P�����*'�e<y��rO��V����%Ys��6�M����^U�QR����&�lb�H�=�Rxg/��������#�8�䭡8�'�!��-~s���>�֪ڬ��8U���#1�e&�1?@��s!�]P3��<�7t�������y}}m�����:ܷ~X�mj�I`��D�h��0�D;R봜lK�G�*f�?RD������D�����,?k�U��"�sv�5�D�M��aQ��~O�d�D��Ȭw 9�1�K�wR��Є��+���s��2@M�;�^ee��ċ�n	����A��r��vVJh?k8���C7�5���b��t�\k> ��l8�ΉE/0{�ß,�}5�06��o�y��|4�SVy�����3rtH���N�b�Y�y�<�K������B��1�θ{��yfP`��4���A(��.�0�r��'	����f���w���v��y��U0�m��X+ ���	pk6Q���a���Z��F�Bد���ΎIn��G���v��n��<>/q���T[���P�I��)�a�IIuxa8%"�w���{�I�D��CT���I��Yyrz�}�������u���gg��"��[G�^X� �J���>��1��+�ԃk~����:�D��B.�ߏ$����b��Y�rP]����x��R`Gl�;� 2ׯ����=���I����%[�-�B!T,6�,����u��L|��6�6;�W�~�[8R1�v����T�Z�+��sc1�v�ط簹"I�:�Di���ͧڃ�"֧�j���U�0���6��-�=��`��j߱/8�Ş�s��徔�$����Ʉr(\���n��GA(p<�I������7����D��M��kb�d�*��?�_s� ��h�=/��\U{�gz��q���ïN'�ח���ΐA�����'���8�W�0d��4�^��$�'���a���/K$���k�Z��U+�-���<g���^��@"�do�|Z���5��o���VyIg�̛V��Pݘ����k���"]��E�j�G�F��CVˣ1���V�>J��\���(Y�d���B���S�O���?
�U��Fi/������w���Þsy�:ɡg��VW'�\R��xK�z�̜��[���5޶D��^��+�u�&�R���l����'s�k2Ύ��%�>���� ?Tf
]�ɳg��.��Ҍ�e���=Xո����8�ڙ��P5{� �b����J�<�]x���?�|`�o�V>q^��ǅ?(��Z���E�<R�������1�M�ɑ���
���j�)/�e�#.�/����P+qѬ�s�tq 25� �1s�D�Er�I�rF9������ ṅ	c�-��N�`=	��X�kءLR��n��^շ �I��Օ�<�������x�AX�������4/�1C��� �1<<��g� �6/�}�i��u�ڨ���b�5��K��9���NBJ[1 ,d�LV����8�G�k�_��_�����E��GC���~<ao�#��a�;�o�5[��ݒV�婹�g���1��ƫh��X�����瀽����06w4U����8f�$m��Tp�>������W�b ޢM������D�n[E�R�����<G��5�P���HF|�������� �a�L���j.�fl�*n�lZ�h�C�R�*�,e�]���&�lZp�?r\t�ǰ9��*W5�e~�}ns��t�=T��c��T��X�[m������n��J��;��& �|�2�	Wj�����{�z���ҜEx��j���s���:���~H���M���y�#���A��>N��;�jVz�{K�A����
Eu�s�!2�34�!����U� �7�"�K-��i���A�X�b�X�JFN�YJ~5��#4u�'�_�c�D�u#���u�w���&��$>X�P J���g�[ L��_�\a��d��rt�*�����B �ei<��҆�8�7�Ty5�J��7�Z�1D�i��F@$�0d�d��P7R�Χ5R�DG���u��fkQ���(���D�M}�%K�2�N!��	0%m�h����K�`�ɛ��� �}�܍��V��W�oMrs'4fB*����~N����p	� fZ!r�c����~�B3<>f�f�'+-+��ܔ�ց`�`6������,���� "��%�Yd��AZw��pg[�e�ii9���(��b�g>�_��7�E�C{�-v�EEM��n7h�6?���@e��b#v��h�~n�2b���2*,1bCӯD�)�^�ŘK�9#ʉ͙�J����g�1�Gha� uZ�;@�Kpq���Y�cftĎ.�ϓ�Y���	��c��^A݅���>q��r#ng�5�o�ү^Ь�dI�w��ڳj%���Ġ����h4���v>>�"^���*.�8�p�Y6�E�՘��y������@=Y�׷TQs�c��?�~H�V�d��?�Np�>���u�������/����~?��$�Hy\;�Z���l�K�d�w�{����@5�U0MxgX[��>f�B.�M9��$D�p��������gQLB��!~����?Y�%���1Ρ�������ݖɅ{�EnGB�i�қ$�x���G:�p$� �"`ҋ����@К��bH�i}}�o�*�:3.#���組|�q��,���e-i!9��p��JK�>�ؓ��l�����P>
T�
�I�����0de��y~-˃�����_��u:R���5�S5+���#���:�J#EX���l�q�U^��2�.$\���h]��BS��1��X[�cb��X��` @*�l�����0Y�e�����|BW���0�iT��y�V��bXu���;1�%'X\[;�	�19+7�7Z]�����������!������1���}��c˦yiE�Q��L02h2��%�PQ�tG��'r��K+��]�^܏�[bJ�eT'k��Ѷ�t�_#��Y:f���P�@v:��p)a�Y����$M4�����!�Zx!1Cs�X*k�(r��k�{ ��V�Ð\���'�,Ɩg,�����!\}]a�ᚏ�D�����X�������a���{6i�^��:ǉ|���#^!�{������E8Kc�~/W�7� 2\��VR�Ɂ�AɝIne�M�����2{�u㋭�K�'�{R�
�gۇE�#rkg 4msi��B٥�������츾��2=�Ǌ��A�v���
U�5H�3g_�Q��[徳P%�Ҵ�DW��Q�?0(���M�1�԰���b�Iw���P�x��(msG�v<��;�mlL�)����w�PF��H�r����g�:c���]�g�t�T�ES.�l䍎����Ue�Z���
u�O��	܀�u� k��2�@(��Y��:P���������:q"-E���/ݰ�aE��|�V����T���a�2	�͑ǎf8�ڹ�v �6;U�rc�Z��}�W��V;�Aω�N"tbl�O���D�Cc��I���+^�"h��O}N�t:)�?�/��%3�`F�;/��l_�y������F2�ۡ,�n�Ƣꛑ���D������k��Ǔ�`�o�o>x�`M����4�7M�b=����B��pԝ�C����X��l�����P��rL7U�(���=�ųߜ�51�����)t'�Þ{cЃ�MA��RS�Q�q�}�f׫!s�0?��M�h��7�I�MS9����}��s��#���ޙ-���R�'BL�T{$���14Q~���
����[τ[Mu��V�\T��'*R�*&f��K�-��p�D�ؖ��%��
9w���L�Fw0�k0����'��� -qN"_�;���l�Md�)DI�W�o)�+���n֐_�O�t������3����=
�� 0�kԸk�)�$[*����ΓU�f�7��hnwD�P W�s�2\o/�4���?;��?�<?f����C
=��9�V�u�[FN :@�5��T�a%�h�����"\荪�
�˂s*��_�,<������m���S��7yӿ9��� �����A����3�]j�k�֨�tj���פk�,4?�aMr�9���,!� ,��޳׹���@��j��?�J8��Ѓ��8; ��q/ك9u�Lm,x�d�;B��q0������C��Y�{'��{�	�j7�vlN�}��z��c*X
�7��ɨὪ��n̥�L�s�Gh?i�h����6r�����wȂ��Q�K�N��'���ϸ�񹮠� v&���6��Tb����ek+�7h!C��rˀ��(v���vž#��a��cM�D}�J/�-}�2F!�w%KF����Y�T��[�fX�aף�/>^�c���Rz��.#���AE�/��+�E6qh�cf?�q����Ŋ�R��s��)�����XsE
�.���J���	�z�D$c��>r�_�4a�܆*�80�`W��m3��&'���z~O����n��T,,=s;<KX� �0��i��Iڮ��faY��8�8TV��%N��6�ʘ��T{�d�u��Ī�C/��X����1F�e�F�P��5C�:7�Ճ�a���^�p�\��a�e�悑t�
�-*���[���!����ݵ
K��u�to$�D��[ �0R\
3��t�`4��?x�U9��i�V;+�糮P�i mt���/��z唖C�4E/y�Y����=�P�D(����7���� �a@`-"ɦcQ#���Q�9;A�ٱ�)�^w?!�(φ��͇ox#�9�ZBP���H�r��K �c4(C�c���Y2��_���Zhmw�q����$�ա�O��Mi���0�H��ǃ���-ܞ/ԩU�?ѵݸ��>���Yt�w9+��>��p
=�k)p=$(H��O�O�X/3�i�>��p��*�R����zmk�*Bz�Eţ�0��M�,}6`�4/|JKAj5�#\�-�^� p@p�"�ޞdC�4���@V"П�Z~��N�d��?�g�[�4w�g�~QR6��ďE�_����g8ǈv�^�llW���\ 0��^q�;^$� ��#*\��
�A
���R�p|�4C/�$�9��'M�9��M�5(ٮ=~>[���nu�A�L�+��	a|N�BV�3m��I�5T9���0���~%�+(��UN�6%z7B�F{odf��6�1��zK�~,�pgP���FT�>s9<�giN�<c�yq�a{�"SK	���̅��s�W�l�u�J���_�V�61V�A �g6Iv#c��D�������������*��c�!�b�̻��(������;�t�������Wp�o�#0mȢ�y� l��6��d��������HK��-$Sr�U��vMd� �j��a�#ط������Yw�rv����UR��E�_�GXV�NEP �����R|ݪ�9����}��q ��Dv�V큥�(�ͮ.��R�z����5f���
�Y���g-����7g{"f�¿�P���9UcyՉ^��m��wRC���:�+�g�$Y䈈3��79���%|��PM��uR�}�hcXQ�������yD�u�NFmE��W��</�{��̳��,a٣7��L�k��W�S]���A���\��1f3��(*U��O�DB�1Z5��:-!G� ?]U�h������d��7�~����e�����~E�����c�=_�.DK/g��L���f�B��[��B�wJ�E}�|�|��\č���	����bc�i�>��o��t4���|tn��9畀d�BT��A8WQre� ]�^9�R�7s��f��<.&�u�&�w�,ԱT�8c���>N>�yRT�d�V�ûA�Y��hr�_����WO���/���F��s�!`��X�2$]��&6
�a�ވ��X(Qn(h�S��KI։2xx.$�T��;�p�I�M��B/5?wt�(PQ����ܶ}�8�(O{X��N ����U�ܻ�@ӖR�3�2����%)��.H������i�����iZ[Z\��ä>L�Ę�\x:�nB갫=�m�b�w� �����~�	����o��P̎���G"G��������ͯJ�k��v�ܔ�nG�o���6Pha�	�rY�h1��)��#�Ŋ�Ex^�P61J-��ʗ�`?�X���j���J�-%
93���w�q��P����;��Y�VVΦ˻̩L�UХ�q���d�!��ޅ�E����"��!	������ S��v��g*&R[�=���1��FX�s)���HE�2e��̴v�r�:���!�@�(�*����-�`pA�Er�Yٿ��D9���/�$>h�~�D:�d�INH�o�8���_�ʀV������y���¤��˱f����tC�����|�D{����l��r����3�Ͽ(�A���8��WAL��αP|(j�|W��DMjt`E���:P�|�Ei�ν����ʢ�[�����qn�Ί���X#�B����6��k�9����# ��0���ު!��C<�5�ʛ!i��T����'xX�/h3��!��4<OzSh�/�ʴ鰉�ΒwS��0�Z�O�ߏe5�ԀG�\#��зQ՚j�4%��C:e�%�$��4���L�nBH}3=|APh�	@�X9
�_��ƕu�D8��<�e&�%\t>�J������XQ&� �>9Y�@��(o�"A�A޾��=!���ɳ')ع��w��a+_@�9y�*LC��
g��	o�]A@5X�,#�Cԝ��5�%[)iӫ��_��Z�'�C���x�<�n��]2E\ǌ�{K��B9vI�LQ�b����rC�k����t�?�\�"�{����Cj�E>6�V�f �?$\����mJ��|(L������qNo����.p^��X��!��D,˭��]69Bn�����}�xsX�����у�[�x�p���A�=�cݥ���O��-b�¼x,ǒ7hL8�B�b�D�6<��q(�҄S����!�?W�6�kA�`��MF�2��t�{�F�25Րz�T�zpꇣ�2��PL�og�#P���Ӹ����O�99�3׷ܻ��mjnO~=��lE�YC��>`<�K4\����$L8��ÕDӽ�H���@��	��䃁W�C8L���f؂�u,w�41��,'�,�g��%t�m7|��B��� �^+>g�_U~VQ��!a͕�Z���)��|2��=Ƿ��6*f��%�b�;5:Nk>+>���_6=�����N�4T |��Q���o�f3��[�f���(%��	W�*�3�jt��~�o�X�^k�Vߑ=�,TU��pϜ;�J��l�0!�8�C�!8$aIsU�f�Q7-|��I,肈v����gYs"�.����!��)J�{g���mG��X.x��%M��}Un�KQ�f ���Sȼ,�2\R	w��${�8����8��P�=s^����y�YfE`Jf��� \�l��6y��r_e\��9)��=-YM�*'���@t��o�?�;*ؓ'\���:������)zM���9�/�
)����Y��p�@����|��J��@h��4"�6�P�����j]�ʩk ��X_ě�}��_�J �;3�z�ݘN0�h��	OfW�X���sSړ=�/j������؆��$���<���*�h��f�Gᮂ�X�����d����{i��<SnW��g\ge�,u�h�`���Wl�s�d�=:�v5��1m�t�_ �d/e!(jU��av�YlV��ԅ��19��q�_��U]z�f}Me����z{I�F*�p��*�G&/��)�o����ⱂ��%��P��\Zh�eO^�!kq@
s.)�&�Mt��q����GD]�&�e~�R��kt�R5�B�zl����o4s��Sm�
�\+!I�U���_�Q��T��գ��b����Q��	V�2B��j8	�a�m�\z����%<l���H9��+Ħr�ꯘ����Y^0V�d��ח��d�$�%�wq�Q5�'�F<�e����JT�$O����]���Y�V	�i:H0K�^�iz��&����obMZ%c�u%�-��D\�>0��kGV��qdXH�kcy̛��CTU'C���$��R�In����`+$�O��2緑��$���h"�.��"]����
�Z`�a5�Y��!g��N�>��u����%�o�����dQ{�Y�V���
{(>��l1I�9
WM�U�B�­tM�R�sY�t˥�y�D� ��}yp29x���c��E�X~X:��b��5��n�{K�՝�]�ැ�cy�4[ɣ�r��՘#ET��Lߋ�ޤ�	�io���!;�nL�+S1��F�(�:�uc�ᐪe�p�(�{�h�|c�Fw\�a>��nǚ�X��h-�Z'.+�p���˿�6� ���O(W']-cmByف��˭�Z_�c	�h�ypw<c:JA�@F��۪�q`Q�N�p59Yz /��3y�qC�g��
p]uL�j��2>�P��4�#K�F4�q�\=1mHG�R����AV17!kx�?u��N��J8ה�G6��1I4�lN�x�	��3	7x��o��	�8�E��ڥ�r�o
�#=�.�_��?<���lu�Q��;eb{�Ɗ'q<��,�p��'qo|�����_����b=P.I�}�cx��&d�`ㆌK&U�4�#r>��� �?������t�����$&C=���}���PE%/^���~�K�4b�!����ͪ�r7������ʍ/�Z!�r��=2��q��V�L��э��%�����H<u�,��W�R���jj���~ѥ}�	dc����c?�i��F�1t 3�l���Ϸ��J�fp{v,�lO�*�7�
�t�/��Pg��� N�	SK]n�H�T������"}���U��z-m~~O��[ACf�!�C1y�$���?%;H$Ӄ6�N�C+z�c?����vu^��1�U�W�"gl�l������+��y]�z^����x���K_���w�9�;T�wx���m���e��j����&�U(d�[�G�L���f��;�bV}�>��Q�+�K�t��N�M �Lw2ۼ"}�h��҉u�}	��2��f\O L\[b�뱗�/E`�4?=�GP�h��(y�;�k~���������\�ٗ$޷tc�V��:��20��m����\N�tI��e�]���|@@(Co��*A�r.RVͤ����<Q��5���8�g0FN���)�ʻ��F����]/����S+��.Nh:�
BR]/-�&v���4�K��3���Is:�0��ouRK��@�I�,��,��r��"�����Q,���񧹸t�7M4�ڙ;�?R��+��m�{�Dw=U�ԋ}�Ϳxa��Q!!03����M�v��mJ_�ᛒQ$��.�ae��-S��N�R�[��X+�H$S��uI�d3z���1�W͎�g3����t�vb��K3[�b��J�PB�:��R���<VJ��^�-�j؏GcR6���RZ�g��U��^�C u��#.	��)S�J*О�>m�9&�HE�%,zk�(Z�`ŵ�]�K�S:�<�\�V�y75cx�y:��;L?���g1u��rP.!�X�.��^f?P�ceݨUlf�k��G=g\Xl����1�k!��t�N��׊%Iñ<qpt���.�Z�O�Qn����[c�1���ZB�BZ�i	o����;�&_+�0Y�
���Q1(�q�H��Xs=�]�� @����D�R/6�Y(X�$�dm˺���%?X���ON^&�'��lڲI4>�*�NJ$⋯�<��KZ*<j���!�W3��(��_��� �!��Jk��Y"Ì�4�z����3�������;�j��q�HO:���
@�Z�GN�d
?�WO�?!�����ޯW�yB�.Ș�~Y`��|JZ����G�n���WaFѰS+��s�I��f$<�-����U���]�?|	�;T��
�ǂ��a��\� �ҹ� @0$ou�#��q� � ���6dZw!V�Ӟ
��M�8�O/�\����h�|=�\0��ĭ��ҋ;s0�����?��+[��Z�2��~�N^�&���~���{��� =ɦ��Rz�%�|f����gÆB=п	����F0|s��>�m�D�e_~F�Z��č���]G�E�J��Qκzkއ;��n-�X�}��Ee-=�o�N���M�I����/^M9��:޿'~��YZ���֡��6����M�����̲
�L�9��k�2qw(ᜤ�y��y~��$))�D�Je��%�Y	ʸ�lQ��@˙G�ޑr� ��+�Q�7!{R|+�0�Q��E[L�&
ۊQ�S�vkI��ng��>���f��mn����ѣ��H]�M:]5rM�h�*�b�������	�$�Z������<A�k8p��$Z�����nÈ���y��{����L4���3Q��X�-H���:CiF�~��e9f=Mɼ��N�\�%M*sED� ��l1��CM�~��\��?�$�*:aO��bp#K~
b�U9�ue~����.ܴ~*�U;ws��������������T.���J�b���=���?Ԙ�v��Nu{ ƺ��w�+n�}���Ơ�>:�� ��ky!Ӊ�,��ň��A�q�ڤ�U�ٹ�n٪9��(���ga�H�=	]Jc%���G܀�`VO�M�Y!�ȄT�%���ȏ�c�zb��?��-�� {�,�� 
�{��-$y���)G�TX���p���N�U�UE��|L��'`"�@ȑ�Xܘ�6�u�_�1/i��_u�5��̣���ٗ'��f��E����~��-{j��Z/�@�����{c�����_
�wLm^3�F���R_�h�1��ϫ�P��S�/�l�+C�i�s��vB��j'��	*0��?��-�`��3d��L�t�!�e���)�IlTg��I�o��!�(����Bcu��" �7�l�a�*I�a�c*I d��Xkc�H{I#���������О����=Wϻt��A��aT�mmV˰�{c����m�~���~�v�&��^W�˫����%c�o�G�k/�4Aq�z�܆�U���TQ�3��~Yh���&��ޡ��HE�<� �b�����U_���\H�+��u
���ӱ�p�m[Q^))�d�g��D���7C��R��.Vخ�,�FaӪ�	o�;����UE7��>~l��F�]ێ�k�cB6��-�tǥ(��u���O524)���/�3F���[���T
L�5{�{R�g�\.��qot3�MW���?�����t���e�34��DdJ"���5����#�sC��%�p)5�^b��^x�mC��v^��M���}�Y�A,����Ab�[��lPA�����g/g����e�P~���q_5#��I�G��t	���|Y	�R���m8p��>�}�U:H$6�M��f`4�LnA�ެ�����]��/��w{.��`���9��u4���}!0�f��W���W�C_���c���۟��� ��,��W)��F��a��A��C��rK.��Q[k��QK%��gL-��ЀsK*%�H"��P���ݴ��B���+����_�9��a��0�h����m��cu�J>���]!�O�g2�P��N]�SJ1�Ҟ�!����9������C�ۄ�T��Z���|O^ t�ϓ�G(0A*�v�D^��|Γp&�y�7�m>
8 �zG0���6����\���o>���ʋZN�S�>_�נQ�"���z��,�w����]:'g�jMqG�ω-Ԅ�6 \|�)���Iw\H�dZѹe�iW+[�y�_�٢*$�
C=�(S�X�cKF���!�)��|RլْU_L���
��ʊ=�N	�'-L9>oJY���/@:M۬�sݸw�V���eC����9�3?�g�P�i?Τ�|8 ȁ��Uth�>�=U*��wg��ڝ�����À��ܵ��ɨs-�	Z���N��]H�׷�n���܈��7��]�e*������qH�/�C�H/Ӭ��K�ήf'��"Y�L,�϶���1� ���k)��>��5���2�q&�&��w#��f��v�D���'�Hd���Ș���2j��u����Q����	C0�NSǈ�=6�Y��ӯN��#
���H#`�1��6:3��y]�dj`A��O֠���DЯm�(�/�?Ɏ��Al��@��c-`��"R����ȋ��;�,� 5�&�mˇFH;5���=�K��@�����T^ԛ�;�L7_�T�9p��$����S"ރ�	��_�s n��9M��\R6	���L��F����Э��rC�I�lh�_h�ο�[���W��#1V3��R�wɭ��@J�#�
����z*OTx�3E�����|ˁ��ư���~�7t����_�1"
%QVh�ՅQ:&g�Pj�uH���1�_3c-<�,��b��D��gȂl��D�ک� ���?��@�kW�6��8�)%r���؅��D��5X�C~�A5�&��v=�����ROjH�YL�?_��8?�\R�I�,�~������C`�JX��ӐRǙ��#���ҋ!��zS1�Q�*�0�j��Z�`��_�?ҕYB��l���E�?�F��@.)�I��i�v��ckb[��;с������h༽����A{���H��9}LTG�"��xj�e�W@#�S%/���eG�C��#͛��y��=O!���2��!���"�C�x�pDHś^�h,�F�I�I	��>�<�'���T���ȯJ�%,�q�7�5;�4X�6`F��A"�i^�k-,<��g���H߽�_��\i�I��*��+����[y
q�����-'���\��ҳj$� {�vNσj���}Hfp��t-2YD[Jɕ����B�g�H:N�%�--��Y�x���_�G��`��*���e'ycBǡ,�)O���B�� ������斴�V��xӦe[O͠ܤ ��֋r�@Y�}�_��0/��k9r̤��Y�Z��1��K���ILw?�$M�9�I�"ʩ�(]��o+��ͭ�Κ~Ti�=b�_m̠x2܀���(0X���J��<�����^?`v�}� � �(B�`�bg4&sE��Mc/���F��?"�}nP���aw��;�m9ᗣ�oO�&����e�Y#�ߎ���<�5�����V��Pq���U{L�
�y�;��3T{/�fC�+?}�:
7���G7m���qB�NLrg�Q�O9>,Q��N��x�`=����-��Gt�鸅0C���Z�uR���0�q��GWZe��*TO�3`C���5k��E�\�A�,q�E0ʌؾ����?���붣w�h$8/�RE�����̿qU��[$�e�1��e�5L���B��3D��X�ߡ�e]xS��oT�I���Ӵ϶Qv*MX�Y� �"�h���=Z�J��O�7�j���ZH����#��a��[����MQ=Y�}�������$���qy(Q�}��vD�ĐE���Ǜ1YGq��m��/&?Nض�p�<�G���~�acrR�up{���M��g��ĩVE��
�Q2�	�ln�)z�z�])�v�������ֈ|�i�įU�9u�s �����8,��V�S7��'M&���]����-g�q[�q:3��3���g����ae���Q�Ί%�t.�S��z����|)�.�9?�6�N�|b�n�K�1�S�#�E\�O_�}�d6���1b�F����� !�X�-�<��1�v`�\Wy���u.7
%�؊�Y��_#(y�سE_�0*:Ftg#:p���f����*8��	R�VW��ϼ�i��a���8}T���y(��\j|�]�� �`��%{ሥ�u� �?�j�"�z�	�nk�Y_hvHf3�r������]/H�S@G���N�EzJ���m�j@3���=D�ݕA�9ȉ*ݚ����lj2$$KR�a~ �2�%�r-�b�$c��	��?thf�-�v�K:R�^�ȿ���%X�@\�@��M&�;2&1�U�O(eƃbA�hf~���������I���qt�-�&B��1fZw�5H�2���Z��UŮYTҔo8\�������hV�0�B6�IW��M�#c.�j�����+Zw�E�� xpԪTd+�)�}
�X,D�5�����%�хP�Hĵ��>OG�ޘ0�o�O�R�T+\uwI����c68�z����Xw�C����^�c�f��%sc�);��O� CC�qz&�zt-Lis�(=�-#}�jrяh�H�����M��z#��M����S�#��uE�)>?� p��QI���?P����t�$�A�P�oV�͛%���SNEf���.#~h �!�(-�5H<���\��6ch���'�B��o**y}P��?�Aǜ�3�J[6���q�t���)"C�~���4ۊag�u��t�6�H�s���?I�s��BY%� f�i��5,���9Yږ%S�Y/�����e����+�f��r#c��Y]I�9n>w.�è���	.���qiGS"�{tٵZ�ʋY�2�̣9AǶ�!�I�|�1+��}ԟ�A���s3d�y肷�n�q,ē��ܚiQ�{D�$���Bv\�Z#
�ibH *ɠ=�$e`���X�&��*��}&U����3�6P2$��1["�U�a��c1��;:��s�+Sn����Jv���^g��*��0?�P� ��hڂq�Q"]�����g�����j���;w����I2@���ʮʗ{�g_�G���>��q��a�v����؃$4S���*w���e�ϸg�]9�ϨGg_��G�X��ש�_Y�qy�B{VӲ7Ͱs���w��5���zs�� ���6Ic�Ԅ�"�<�z\?�|�����x�'�l;ܑЙ�ǸG܎��#Ӷ�ҫ�J4�����#W�^�v!YE?A@�E-x�Ϗi/<Gm�~f �v����(�n1E"Kj̀ms��2����:�٥Ђ'����W���*�Rb��.`~ju��|�IO�� ۆ �DD(p���Z�g��^�'�8��#T��2j��MpS���4�V#5(7|)wd��t��g,�<N��A(��lmV��$�,v7��,�lo �˴+��^�~o� V�j��S�Y�s��$gܾ��A~y�X�k+���@�]^�����,~kJ��l����JjT(� �*LU�{nA_�����H^���~ՊwW�/"��8�ĬA�D�$��X��� �01 ՞V�����0~{��]}tC��Y	�b��U�ڨF�{+�/���엞$��\0��>�%�p�ɂ ���Y��0�~o.%� ���i|
s����nXj�(JO���hbo�{��eh����uf<j�t��w��ۤ�?*�����cd>���پ&��QA����>�"���9�o�@n�nhu�b�L����^2��6�����z��V`B�e
���W�v���FY�7�߬�c��n�r�o�FO�Qz<�z�Anʅ�NpY6�aY��ɞ»A��zi���� �<�1{E n���N����^y��}���#/�2��Ef db?e�ż@���S�'�b�wd�ҊՇ3��Fj���ŭe�!E��_�f�^����d��4�)���y����ax}�b���)�6=��:Ɍ��-�P��d�wG��^ɭ�)���� Y� ta�|�v�<A��u�9F��$j�В\l�j��8R���NĩK:��Dv�Y��sL���3�N��?�+5P��  A�Ia#�T�Qc`��v9U"_��xCA�LΧ9
3q��F�Q�_\�bɂ=�(F�K��>8Q��`-�/#(!�C����3��#@�^Q �la'�����&�j����ܒ��f!3uN��st��W�.�3_�*�?:�Zʟ{F�= ���+S��:�V�H�����2nbU��V���|�ǹr�|�Fc����X�rXRmy�/�FT��'�+=q-�Å��I�"#�7낵b}BFWt��D*>�����*ap�欎`H#37�:r��������~�Ȏo ��g�Yaw3Z�`���*�2F +�Y�݂��C]���U*� ����G{�[�紀iスs�3,T"�>�H�M�^��6{�}�]���")���x(`�R���..�ͬ#U�w�6���BQ�avs�{�%�Xw^��4��/�
6�;�h>߈�\�����-7�@;5Z�-�n|��d��0�J����Q�+���R'��$Q���B
�-�{A��'�{��]�X��c�K�dX�?��V�Y)�n�"���DΡ�c*���]{����[ՄPk��H� `Aҗ������:����d��*�7�y�k?:�����u�)�V2Pu�=��i�58KB��DUʋR��a<�J:�3Nؙ�������J��2 �Ug����9�$Y2�v�m�SP-���.�xB�7,�� @h�G�n$�yv���-�8��8���e�͉�&g��虝��܆(P�$/ui�رl��7:�5��=�#��X���U\����rN7^g�>Jq�ð�M-��35c�\o�����4ZW&�rG�k/)m`��o��u��1���*�>�o"��s�M��-&D�ȭ�P`Ӣi�V�$G�}��)N%C35�x�0��lv��C��u_*�ӻ1���g��~���3*\2ex��5�ڍpXמ�u��^x$��ռ_	�?�#�����
	�#�P��A����)�ؿ	�x��i���.�ؘg�:d��·��R�,��)��;	����P���,�y2pNX:�jz~��S��GB��6�I��r����aӘC�_vh7	�D�w�E���cA�o=�V��$����n��Ƅ��ゟ@��8{2��t�j��L .����BS�!a���<HٚFYI�7�!U.q�ai� �_�BMR����+�x^��6K�*�Dei�����Vt������'KK��6{�·����TOV���'��ؒ�<��EStm9{c�f�w(�	�v٦�d��H��H��M��Lp�%�h��0U��'cҌ��9~Z�8Z�k��4��|�����I�"#����Z�<��2��Y��g���(������G�M[0x����@�̅z?O����aF+�?�L��}y��'�{�/�fz_���_]�W�v�M)��A.�T�e:M�O������ɻ��%�H����ֽ*���|�y��@�b"B�����o����p�CكqC��SBSwЕ��J9+��z�&	���(a�����٨q�#Qc��6m{��2Ճ[e���͒�(���|,�^�=S�0Z�� �51D�{�x��1���@ɮؙ�%/~h��/r�_�)�8���|���Ɋ���	h�5�ɘ�0���m�d�`���X	��E&$�J-��o	�Oß��"�a��w�.g4顺E�H��M����Z/���Wv�&B�p���$à�q��S���Ň"�؆t}RU�U���=�t�<�e����4���+�)N|z��g�#�9�%�2˛Z8��� �q6,&i;�
��'E���~q7d� :�p�=�8���/Ǔ�A�u^�|��9kb��*�V@Y.�"|�% ���)��t��<���uq 4@RW���J��X6��S�J��a?)��r'١g�m�mOwH��39�I���{��7�<B�'Z!����YHL>�� J\:+Ϛ~o�Ci�膭c��'�c�d�+���	a��+����$���]�S+�NU��*AY��F���K2��������O���Pm����kt�85�l��	;�]&�t�+Y����:�Z �R�|Ƣ�ڂnZ�d�V,���3�>}9V�2��o�d9t#���� �[���}���ﾗ�(ZQ�^OH�`��g_*Ұ�w95�]�.
�J�C�5c�v_�f�D��xc��M:=}}ႊ�T�5�xP�$�?e9o�7�AÊ!�"	c���37Ɯe��o�{Hi�����O~�9����S�w�Y�����9L� b����@�4T{�������dX�y����${�,Į�5�	��fB��z�n�T�0n�@��48G��XV�R��UT���6c��4�$.W!�1�{�Ib�b������۲������� ��l@�ۢ���%!�=
3��A�'�w5E_Ҋ���)��$�	ͥ���xg��~
������6��+�*����Q�M&�~ �d�h�:�����nV�<йdV�<)v�_�O/��r���~o�hw�Նnl����7���p�}5O�OI(��dv��d�RzV��Xd�L٨�a)T�3qm[���|a��<}I3���5-Wo��BXHE��|�`�k޲�N�*y��0�f��_�Q+���6V�f�I.*��1n�zZ�0d�7@U@�^��]�,+-w�<=� K焍t0�-��ci��To�&�B�&Ǎ��$Ew�� �Ŧcc�<W�sĬδ���>�ߓ�(�eL��a�%nݎe,�*8~Y��=��%�^+Dz}�`�v���>��lMcT���dȨ-<�/2�ܐ�ذ{�.W�'�ȓ�|�j%L�c��$����g/�!!!(7� ����"����09a�ϲ��b�������{�.�*!\4jS����xO�!>ez&��m5.����o��{e�xu��|HX�8n
������#IIS�7�~š�}S�%�ma��������ZT��C� �^x��}uWHq��l:U�f��21�I��<��b�?a�6���4p��X�����5u�U�B3�	������Fl>>�d����7�]���2=�F��	�D<SeV��?��%�Q͚�,2���� Qܣ�[B��M}��"�S�&�~���NC%q�(�l����\�f��6M��1�ܬiv�GU"5N;s�2/�K��\ֱ��=�݆~�8��rX��4�mw�9�T�Ԅ2�a�㶒�щ�k,A���ݬiG�V7��hU��=��t��51�����]ϥO��E\�2� �̀@` �;C�,QM�U�|�K���{�F����Lz�|����w�*b�F%�é�M}����(�fp�9X��O�������_���M~�:˼�_���8�]K:!�
���F�%�@��{�)0+hv���a�>h��!�:��_��Hz,��ܠwl����<�K=YG%xf�oP��N��.�MO��J8�^���z*�,O��d��5tV��JV�ô�R��s��� 5�H�_��0��[Tw������6������]p	5r��+�v�Q`����}�IY���Jg��}��H9	���(�@0d`3�,vA�Y�G�yHr
W����4�E��j�e&�6/7�|U��K�WW�`����2p�����k���:Q"a�C�p>/Vs�e���b,q�ב���u�t(�(Ȫ�ֿ�	2ʯ��%��:��lvh��Z`s���咹Z��~�Y����~PE�-�7L�/y�S��VȆ9�p��rMV�)���˭m�K�ݮ�s*�.�#h�2+9����DK�����5����M(�	
�ꦵ(�(��m�x���Ȃ\�w��d������Ogt���}w����$�bwL�g�9A�0��FX�.M�P>pM�Br�$X�L�$e�F?Z���[�c�d�t���o�\���� �4��h��9��9�%���	e��ݯ�r{N}<�%J�uߚ�;���Qa�ے��N�O��`�u�l�;b���e�c6�����߼\<>�K�����=>)���D%�w�+ͤk��n'F�;*�`6zt"�ϲM����[?qєo���qp�¹^�b2�>m|�?RNS�g�D!vm�Q�� ��,I�IKSXi�^ܠ�d9v��J�6�!:��/M��^?H�A�Tc����CG�n���d�60B�\h����J=�c��
��>�c�%���L��d��Ѵ �lB3Wg��'T19( Ϛ%�)��E}]�(%�7;�_~'ml�]�k@o^���cZ%^j�K誾���k��zK�#���u���"�̅�
u�r�S���4�^!�~���S�Z&B�k�@�
�M_���'!�4����	d�F�{��2���,��ݹv3w���H�X�aOB!ri��}�W
s����x�b�SYFa�͜��4�ү�Eթ���jٓ,/*����k�������C���'�J��-��?E�1�/s*a�_�j�ں�V�!d_�2tH�������B�k�)�N�җ'Ǎ�������̛)e�O}�Nu��Q�#SM�-�kťg���O��]+�&���0�M#���������Ȼٍ�2�	��2F>�'M�h�uw#���c |� �׃]�uw�n�f�/��塗���o�JniIzT�.尐}�O1�k	��f���$��G�5s�ʦ��:�1vӿ���%�;�k =��e�A�v�#���/���L��!����c���\�3����+��\�	�dYz={�5ni2�y���,R,&Aփ(�ܢEoH�zد�w���$K,�֜��ҍ)��z"�5W�ua�a����׌.$���/��T$D7�Utp�b���$upVt/��������.�ܼ���[4����a+�ed�ڽ�ao��'Η�u�c�:���ÇI��w4~i��؀`�ޖnĺ�%��" !!g��iJ�m�uR����ZUk�����/|,���Q-�􀣈�!?r�Xdf;��Ivaq������L��g���/v[��!z�y%��o�2�G��9�"�0�
����u��~��+s�T���3e����hl�5i�Ԝ�-�6�A�&Л� vT��}iσ5���IJ�SD�S;�*$4�����F��#�⒂�bК̚A�p��F��3��uOkR�����8)�R����ù�p�BQ���F��Km��<N Hl���vA^��b0�ui�-�(!����m4h�:8�5����OQ�M����>��xZ��BO��(�����7-��6���#����C��?_~':�ٿw�?Z��k��9�x��Lغ�Xpd�W��o�d'�������	��嚷�[�*�W�p -%;(�,Et�N#�pM�����nY�a�ͳ�m��LZQZ1J���)�ƈ��Eŏ��k?Fʒ�#�������NQ��|�z�C1k��s-���g=�#��d>�vG�h���Be@�/��5`ؔ
��$8�К�9�v,6�DYq\|#an��5{2��T�HJ+ٙy��G>���p�^�I!��P�a)���'���.ړvK�C���aU��;�#l�����掍���z�f��.���T��Oi��І��@Q������#?��6�?1�7H�5�CZ��g� -����kyi��w�?��� ��?N]�h��l��VU{�۱��3G�C�6��r�P����	�(t�<�n"���`U:���#���?�'��[�g�:`#���:�K�s%.���I4��[WK���h�5���b'd�h���;��׭�`8®V��������>��w���dqR��<���hK�l�Z&�"Jd&W��S�3����$?.�TZ.\,__�e5��$-we�1�e��ŀ|��*B^�hE�K�#Tv
L���^T����o/q&6�$�h>N Q��8��o��]�\�:��_	cJ��:�A�j�}ɿ#�J3�GIuh�@�� `�Ex�sp��V��16kS篧_���
��%��~7�63����A���	ֲ�.���@����W/h�W�4�O�fESؒ����
�a���?A8>��<@���&4�h�D��]3E�3f�6qn��n��g�3���;�;���2E��)�S��
�V�vڣ�T�U6�s�	F���EST�sD�\
Q���>e$	ɫ��@_��\n�e��ݓp��LC�tC3��.9�2�K<��=���/�������l��Jm�KP!�%��9{�eI��-M�vV�g�1��"��ۆ���4����c���ϴ�����)A�Чh��Z��|��O�h$��V,V����S��� jY9��}ӈ;����w�</Umc��r�ް���+����C�tnX)c���n�
njq���
��>�G-���!nV����݆�
�s�Ai��#�}��㱹}3��!⠗���� �\���������լ76v��H��M`�Pg��Dð�H��,�&�R�d��PZ�go�D���Eߵ�x��aD���h��{���<^&�.��~���TD��#RF�ؗk^g��s����D\\�r� ^r����T4�$�tWҔ_�ֲwŋ�Ԍ_]M�G&t"wF��W�œH�A�ՀZG?��Њ���-f*�����A���Mk�H�D`%/5�=��J�LmD��������60��	H��HB�miS5Y��e�6Z��Op����G0����ܕ[>:��\�֖�kD�0��
0'_�4&D��z�sT�~��Ub��B�*� �)����uҒ�c	��Nw� ���$z�|�=�~��OC���<bn*���j��|��0����NUF�Z��a��v�0����wM�~��꾭��w�SsE��>R"���F̚�z���D6���ɺ����V�m)g�ؔ6 ୖ=�6|?���0N6&� ȯ���6g�G��eX�4Kls�su�	x�ͷ��yv�GSi�^��*�����ī�!kfw�NنGg��rߔPE�m�\}܏t.f�3=��rⱔP�^��.��M�O�AR���/n�E�@ަ
zU~��J��1L�G{Z��-����	������~��z. �T50X=͝@4&�P��)P+�z��s���O��<�y�m$�����^˧Y�,Et��?YJȿ����٥z�;��I}�=S���� H��r SaI�����V��P���c��:I<jK�U�	`4�t�Zb�p5"�j�*7yl�-�dWC�8ߏ��������䓄�|f)}�[�c����ټ��n8�ߙJ�!�=��S�e��	h��A�������QZ�K�--#���M�HF3��u�L��n��ҥ8C��|ы�֘&F����Y�H�l��� �?3��a1��I��ݐ��
ݫ�:D`�9{
Z#���ʋ����2��>o1��ѥ�F�9\D\[��9n� m͋��"<�����ï�~w�C�(\�p(4+�����\����0{XDB�,��\PL^a�4i����H�`�3=2��^9�a|���ѹ���#x��:O,[�<kAq���zw7�/�#GN>V�<4��%�7�U9s�� ��oq��v�/�:!L��[*�w\�,�pdkH���P��L\1K��J��	_N~	G�b٥�����%6�b��"M�P��'{U˧�����mω2�e��)g�M���ۆ�6�n��~SwyLز]����B�M�9�d\�����tŃ%�h�kd��2��z��F}v�y��)i,�9�4t�щk	�I:@�.*6`ؑ�CN}O�j`p_"z���:����Q��^����ik�gv��e�5�K��r�A�9����qt�!�]!N�Z�Z%h���i��]�Y���~yd��b`^��>s�ݦ��M��L�5�t�ƿqF�db�7u���p�y8ܸ١t��Qsw4]�rtaC�4��.G@�T.g�����PP�m~7��j5������=j<Qq��0`׆:Nȡ[> +9L�څ'� ��(\e5�r�28D�U8T�(/Z�j�`oh�
G��r��"�]((:��8*��K����D�E	�u�U�X���(����~T6i�E�`�՜�p��b�[-���yl��P�W�$�c;<���EpH��u��r�&����>S�Vp;ڳ#䇤���˙i�\���;V���w;�g��.���a8���g��<w5�j���c�IR�>힚� ��aپc�o�A[�Uq�F�5l���<��,;M$�$~)q�3[��~?��lp���E���ZK�؇��3�ra\e.��4��=���U���ł��V&�,
CJ�M6�\	BA�63Jq�^M|�@��t��N�0�2�Yv�~��d�t��:�����,���F����fe���,N���Z��N;�R6V�q��srM�ēi�XI+�r�#XG렜�e8@ d/��n���\���ÆY���o�#��hX�=�1�`ޫ���u�w�CA��,J��*�yS��}1�6(`&Y���<Bd��������P��!��O���C����r���&���Mݜ���2~�A��>���,ug����@�o�iOL
.���]�M���M�9������b�i:�'�4��������X��96m_����ڋ��E�Oܼ忼�D���WaE*�_K�f_sg���-�t���
�>�*Gy�^��D&��hU�q34ң���&���_ea�Վ���Ŝ4�yh�"5,M��aٽ�{���/��/�nk
C�D���"��0���D�q��)!�3
�aYu���xڽf�[���odȮ7�t�{2���g�t�����Z��dXϫ�+�xfN �h� A:< MJ&�W{��������O%5)�q_���5�ȱ�0m$JҜ�=�_9�J���
��$1t�%tf=Tun���sF�Sj���2�Y�OYs�^�L��6ȳ�/��A%���߸໐�#�knx�h����m_��rw���k����6�%���߉�����7�wœ2�z6EȺȄ ;!p.�Jh ��|�7����,��A�r��ߔ�����%/2%�`L���XU�`��d�ض��|X�Ic�)��,dW�] U͝�:�+e,���w��c����=R<.�J�M�wB��	��1��t�	���>f+F��F FR�5���]N)!����Ž�t����@F�e)�=�j����z�mL�|C�BT_�������#���[p������4��+�\�aZh��H8�?V�Wɷ�,V+�:��ALU����_�~��G�O���Ed�H3�;}�4�z�����5��ߺm'�X��H ����e\�>!��3|TJ��M�����=K �;%'t	��(�q;��-n�W���3�?�%lm�I��u��|,=9R^���T�.�J ל�l3���5@���������˒><g�o{�,�̄FRj�fW��-G���g�;!Y�����T�҆�~�+����n-��ږf�#�'����D�q(��י�f�/�Y�i��҉�b{kםB���O*�7mܟ�3�E�_dRc��`�ؿL�D�������I)���+�;5��*CZ�������g�O#��#|�&��i�{�^����(�P�j\��	���Ȃ��)s���~g�l��'�csY��CinV��CrT��=8Rn�'��u �,�`II"s���%�6G�e���"��i��� ���쎏�,�{�p	��k�wV0�~�t��%鳨d�DN�y��g���6�P(�\�4�4����4�Qqn��_ri�y�Ə.�Nw=���WA2Q�-��Y��N����%�J|�����T�����/^ϼ���s����IC����m�`�n6�������[d�	�w@ڞL�䈪��rj�P=ދ+�՝���*�Cy/Sy��C�ίH���;�nDc7F\v&��4}K\!�/��Y�EM	����@��P)��
��7��v"�D�A��6祿�P<��ly���߷�꥞G�p��m��#z:�`��a/����J(z�Yqxhr�*ӯZ}���Z�'hf|�����>S_6����`M�g������`!��D.����5&�pEt���� �����2ޓ�O�wt����ଠQ���XRQ'��:Hr�*B�a+����ƽ-gybѠ ��{����⭛ ���1�}8HWv�D��X�����,5L���f\6~��*-���T�f�~s��V$�D�W& �,(�M�����[_]��9�zt^
���2�I^�	q[���k#ЖO�
(�Q�Yܭ, %<JjgFb��1;A�����:Z����.R�q՝�����B�@/_b��������DFD¬^e�7&��,n@E�?�'��5������0My)0�v9ћ�\��f��7e�jҴ�o��A|�����%q��yBWE	��{anZ���.���oդt9t�v��޶"9t���1���B�l��Adu	��iD��'��(���K%��_�m��j,u'�J���m0����8����k�9���DzSBsVFԼ�-�W��A��t��?p���5_p��wc�g�ޘa �� �yƪ7,��'�ZxY�l�F�5���';B�d��n/+m����k���u�uױ��WVD��F����S[�9*�ږմ��P5�瞅Q������-ї��K&_��pS�z�O�5��o�dk�t�[9Re���)���<��U8�=J�/�^+�&2�|���6�=vH�Ͽg������<�#��.C�z��pp1�������O��l�57ت��� �����#�2��T�?�¨�M�,�v���w
u�޸���<���h�zMT�;��u�H����p��w����Ǡ[�PD��R�->��sS�Xi�Ѡb��*��{@��x�R��5)��)T�������ђ��������e�����.?�؇s�b�AJ�	���	�v{�*cfΈ˯v'�-���0K��EL/�܋�N����)���|��:���hӎڂ�[����.�بƢ�ZBX�聾)%q"�t�8�1Q-vBq 罠;@K������H�!u���L�l=��	�.�}�Tm�fG^�. O�W���0�`W�'� Ί��5��O����J�5����u�^,�	 _ �̽���R��/n��
�:D1f]y8<	ڢU�k&�ܛK`q�o1̰�j�a��Qžw�~�"k�D�d��c�+�_WJ��)H�WyP�X��3H�v�O��bd�9A_r�P�}�����g���};^9�ήn�q���X~��� ��Z���R,l��S̽���@&.zPۖ���ew���������=��_t��d���4P�T�V�]�)x��M9�縠��ET6�3�����v�^MX�Nt���@�TD���^虼��	}Q~BdU��Wk���ҽ6Qc��O\���T4����;K���c0`�.�ݝħ5"ԓ.�4H ��������v��K�D��y�I�jE��4�	�m��̚=z�8���$~K>cN`�,�=q9��&N�<�n�ui/7av�u��QU�My��H�(IOf���R4vE@t���ޥh�^�Cb}��`c�@�nG���竒Ӎ���M<Њ�`�U��
�"4�Оl��l5#!b/y���LMB\�\�Ue W��VӦ����Cz�(��Cgo��U��B|�D��9�d[a�0]����M�F!�L6t���$h�#��*��"����z8���Cb�#�yu�ۏ��q�&��`˸�EkbTS�N��
���Ri|�+��9{SV����
����2����b)��Ęw
���e������Ӌ�b�^->n7���R1<B���zv5֝���if�L�O-
ڽ�$ O{�����P��&R�D?��f\�ד�ܲ�_�3�&	 �6�<(������ä<\�7T���w�_�_��U�Xj�J듁�N���
����1
�)"s}��>��4��R�^9:b&�)5�'g�&��e��&�����|���.2��xJ���7ţ}U�A;����X#�L������2��_k�«�%<5������z�)����q}���q�9�+^��ü���!>�u�Eܮ�*!$�r#|u��V,2�$�c���ʵ���޽����Y��И�A���m{���e��K]���}^.���s�.�<r��;�{o�>��P�����Ó]��x���0�*���A�v�őmR�3�o�r��|�e]�I��>"*|u���N��x�k�������<�7��Ӝ<yaq���5�G�e�2�>	�z�3��V��k\��(�#=
�U^�3�������ﶣ>[�N��+c~'���y�]J�+Kb垆:m{�i���:��=Ԥ`f\�W�Y��	����s׆�m�MIn*��X���P�k~��������TjX����%3����I�ݸ��}B�;����_g�E-��~�|����5�a�NK���� _G�\�ʝ��SX���>�c��t��#g ��7�Fc���a�!�����L�a�kO܉�DKMθ=���`m��.�)����n�\�ʵ�'�k���O��� gw�1KP"����qbGG�l�qSܤ�c>���4�f|�N�ɼ��-��ʡ��c��~ ]��Z�9<�f&�O�@��AU_.<Ւ�Hڥ�g⭤b������w���:���0kF�5��`ؒ�/4�9��
@�	?�CZ���6�^ d?L
��@��S�TR���9"��iQ^sUi$��v0콫E����Vh{]�:A�����%���z�O�c��V�N�;�Ԅ=O�����)��}���.�FW�l?�%e�� �ۋ)�V#N;��j�g{"��ѭ4L��ix0ʁ�Y�4����.�ݓ�x��a���AV븨>�Қc
iݳ��:�������(�v>V�G���g�%"�Q�V뜠Ǽ�IN�N���,�2�P�e�����!�?��]	��MX[�D��W�5q'��lKL��%b�a������j��3}0͠Z<�m;-��`�[�0�uP��;f�<�ra�L��L�����a"a6�[�+F8g9��r'�$���
h�K�H˕"�w�;��/y�YeF7`"`��*��W:��8[�d�E_���&#G'g�_
*�����`��(++�58�1�nQ	|ء�R��?�fz?�/@?s�&Xa����r��	to�ӗ.Z)�Z���/�Y�eȻ�.�����,K&j��K�~h�� v���A}��"���|m���'���0��͌��m.*�K�cBx�/<�@j& 6פ{[ȴ�E����-C\c:�&(:K}�/�"�>J/�0��tnW7C �d�[r�?4kc�&^��k�XYv̵ǜNu�
c�g�*�_�C?�]�K����_�=|��F?c�m}Ҝ�dFĚ�_u�'�~æ�oca��v̻EIf�%e�����։Ѩ���������t\"G���~��jXp�$�����w��NNee9�f$[��T���� bs*��|�Ʉ��dꎚ?>o��9��u�h�7�gzŋ%z�(�q�t��Rx1��;���I�܉<�x�|�4i�W�-P�&�.1 �M|�ny
t9#3���Y��E��Zh��O����;��:��]O�K�i$;9xN��D�-�,�v��삘E�s����f��^�@�	<�#y�&<t�0�9���v�-��y��|`�^�t�\����xi�8d2��m�wE�����M�sR��z�|�(�ҫ uMw�f@�_x7�`�C%�	1 ��1��5�8H,�>���!������0	!��6Ib�=)�������F��a��;�%�?^~�8��?}�?�������U+ҌH?'#8b��R+KF"w����՚4��}@uG�|];��=x`BF���l�,=��%���( �aio���ޯ���q�hV�>�*�¯>�<�0�h���4O�Q3"���
�3��KD `��A���d�Gm�4�
_h���<�K)�t�e�#@+��S-48.��&1
?�P%x�+WJd�QB3
�����T{�vP�Q��lX��Fv��j�Ԧ��H/Z��� Y��7y
��@}���x�N�ԙ��)�#<	$��}K} �t�y}��̈������X7:��H�w�fi����؆�N$����T��o0�mާ�ρ/��"� ���324����SPΉڕ*���V� \��KC���M�@�e�����B{�\DK�*��q��ɸ���}/��B�,��<'���vC� ��r2�K�Tjn�bK�*�|	���Ǉ&2�2�C�\7���F���������@�{j����8C,I��2B@A���1!��t��h���>6�caB����&�m�8^��1p��j��3�s���4&f�z��D��,xh��AD��$������l�}��ԑ�KF�0�)=)��+'M�V�� �GP��H���Oc\��L�v�-�m\��2��Gƺ�-��P�3��"��s.M�G⎽���R
a.�������[�Ɂ*�z{:ۓ)���<��z�6U���3gF��'�2	vh��i�����)�d�=x���wF�z
|_��D����qc�\Y��(�H�#�o^�����.�����LG��g�t�t>;ĸ������� d�7�U����5
h�<體aAo1)��̟��תc��P3��#Fl��$���D�C�dW��lQʱ��=,��,�i貔$��L����*��!�gy����%�甅�ӗ�)4*�-#���^I�qN�ʴ�|�2����L��|����j������r4�2�<�V�cG����b(n�9����fc%H2õOk/+5�ɺ���jO���B���q�0�pX��A�KH�6��n�X�A`�1��6�KJP��G�~��p?���j9�+��S}k$ɩ�yn�^�T`�:�B-V
�J��HvFb���X�6d9�7+�H�K�<������B�Ǽ�s�V��a5.j�v�1[���o��:��ێ,�P��Czz9����v�5 �M07F"7��755�Q(=O��-bCR.��_�_D��eDJ���W~�ͪ�.ɓ���.sy��˝�k�㊹wm+��Β�i碟/u9��z�B�������D�����u_;����G��M��FX���">���ٴ8��R�+���&Z� �֞�����:ޜ}OZ�����B�%:=3Je�ҳ��>W����@�SP��)�^�`|�0{���fg�]T�6�]�(����C}�rP���~�Zl���Z�B^_�T�c�Z�][3��愴>��Ah������Ί*w#�Ԥ�$���z��)����ɡN����P��S��Yw=�/��� 52b��K�n{ r�H vz�JN���9�V�t��=Ƕ�~w35}�X�.|�k�PVY�}�>�"���?��vP��l�þ���<����"q�o��⁷�9T�o�ʥ�~?��ރY�o-H��!����h�W��dt�\ؘ3q��æ�&��K`im{ �;���j�
~���v�
��g/(�:���%�[`P�y�ۭh��*�,mUT��PnB�LK��Bfk��>��<�=�Ym��o��{ ڶ맄��/1�����hh���0عZYټ�s�R���c[�p�Y �j��
|:x̥0~���Y� jR��'�C��6F��zM1�yD%Bρ&[�NXQ�P}�E�d$�H�̈Z٠���F�_'�Ǣi�h�����\D�%b�(`~E�[�����8�Z�.����;����?���|�����+t�{Dg��t��B�
@�YD��,�����.A9�[#����p-���� �Be��81�=�g��N&gü.?PT m�X�~���U�O=�W���J�d��$Dk�*:�)��\G��P�_8b�-�J�w[2���Eu"�x�� g0%�s�!�tV��W6�!;&]��p����jP�����v����������W�?��qaC����А�qCO�&9����A������K��6��6,�lֵw)����q��)Ё��1����_Wm����W0�ibh~��j!��43	2�j!�&�'����Y\�>��+�r�]Sq����9�?!b���:S��FZ�s=����x!���)�F��U�ŽM��-��?�jN�k�˄D��`Wզ���u�q'�ꊹ2��%�/%�Sx��-o/�mg?Q7��69�Ob�ѝ�v���Z8�^<���1�2���ϙ�#R.|�Ǹ�eÑ��<�� �������!Z�a�(�5}��1���aLX��-fkX��k4������=K�;�BT��x�1�̠1���m�٥���!����b�s��P��>wZ�+�W�%E�(Z埅��|ڰ�yF�q2����*feʪ���v֨"K��Qq=�0����&2 �3�ϕW�v�R�`=��낅��C|���0�S�(�Q��x���q�x98&�&�&hԁ#,���T��H	CҴ��:Jݡ�O�@���@��2��vX�����1'+�r�c�f����������6S�	�'���d 9��r���du��X�h��ܯP��Q?���o�=�'dc��Si�|��<�e�ndT'�d��-v>���]�u�-�o�G����{tN�8`����nt�휔ʹD�&��"?ɗH�ƃ�X;�L|�@bڴEKe�+��"ۋW�n�b��?��Z���|A���N0���\�K�< l���- ���p��My�7�U��6;��I����sN��ԇ��2%�������ٕ�b����i�ȱyǷNC�nh��k��̈́���	��˼p�q��5�h��c;^�<�����}�8���P�0�.�9m�J0٘+am�G6i;�~j�[��
���,+�j�=aՊ`��������]�f%�S��,�2�vU��g`b�B3?�H�X���gI���7E]�I# n�����'�˼n؀�͟:���|���*m7�oѹ���7ƕ8)_H��b&yp$�~3�m����5`�I���v]`�ϩ9[�ѫ��j��q[��c<�_�&���qr�>C��Ӯ�z��6%�T%}-���ЉCFA�h�t�����8ySZ�*Z�)��eX˓u��Я���\�\7�c,{W:d�z�� u���1O�����I�����c(O�B�3}�%�]P�a�Id�(L�W����'i�!�xԿ��XU�QX�`���{�J���4��?�Z5���:oc�
�E6�V6+#ѡ5fW�Jю2�(�,��иf ��/l��M�Bq%I�r�*����rew�
L���^~0���3=�\.�[�y��tad+d'��#.��h"�Q�Go�7�w�(�����=�+�`���p����1�|��xy|=��<��m>Դ�O�~<��i<��k|_S�->��a�N	ix��f-F��z��'5Q$7�����39@d���ѡr�,k�!�dʫ� ����h� ��0͚�K-�YS&�{�~�E�e�*v�P�~�i5��ހ�$��k�t@);9UW=~#?����0RK}�<Y����{+��;�[��Ĭ'���9�>��[��p>zpɭ,��k $D���/�xǹ��������a^��Y�3�����i��S���:.O(a��56���ԫ̼$��rG`���v����a�I
����\��y�`���I���y]�X(�:!����y.o�u$;�­���,�l���o��C��������m�w��"�D\�͸SƊ*WtIp�H�9�w�v�rp��^^��>�u�g� ;���J(�#�zv5�h�	�:���x�SqBt������p���ٽf����w�����k�v9���ߤ�����h&�������A�@� �B�{��"��b)&ێ���$��&	/���vQ&��L5!��d�9�wūD�4�ǒ^�O�rez��bΒ�WL(�Y�=v!�cV��G��ȎK�8�x������e=߁l�ɭ@]�sE	��I�����U�}��U�JkC�:^q�ס��B��q��?��it$i֏��#�N/���9/�t�2�(��c��vr�R%g��D�$ ��8�����Y�E���1B�F��F3��#�������i��x��ѵZ�?c8�����O����%�JI�yX�"��@rQ�B��۸�D�Z=�!���f����BA�D�v༴�l�V���!9H���UC)]ҕ��Ip2
ಊ��|���⹥����7��� v���5�;�5�8.w����uR������-{[����~�>n��˃^W7� S�E+�srw���;���U^�2�@��p:�4w�����<K}�	�q"��B���L�I̒~d6��M���,��j D�E�Y��m1���D��x9��ۧ���]��r.S���e���̺�V���f�c�D:�TP3�V_�I��׶���d�,%�1a�D7�R�5߸�#
E�1G�������D�2��N�V[Z3�4��ߞ����>�B4�n�m��m�	���`
a���^�=���`�J��&j`i��]�ܢ�g (�R��Kɥ��	�	y�l��⾷��gf�7�Qn>EX��v8/�����y��=�!^�ڴ�D�-Y�;�zf���
�$ ����d�Jn�ϙU�S ��Z1�o2�����-�2l�/lU��C����\�e�hsJj��Q�s�D��Uk}�{G�Y��V(�$�0ٲ�;�VMˇ����Y ���~;�K�-R	��Ɠq}��A��B3 �'>�b]G$5��l�"�1�*�F��8|!�z�JBth�[W�:���
���ī��(��VHR`z�a��8دoY��2���a/���ߵ��R��z���A��c/�V�8a(�(��*�7��O.�R�)���,������W�4q�k��N[��t����r�ub|�GHp��<cL$q��-�"��ރ�)ꉊo	�#��'/C"�g-mx�!�Mҙg���v�L�j�]�G�T2��T�.(��8~����JE��	[mm`�a��8�b�;*j���Zfv-����&m��jM*wG���#q,>Ew7Gv~H�-䥂����}�W�<t�N��T��^�%fYֹO��^��:�<�>�"k��0� h����tlX9c�������G�k:Ș��N�(wɸ�vg*/u�x&���|Gǣ��g]�2w���a�`N}��ϟT1#�x��$�^tQl���{�d�Ý�o�L�֙먭:�.��.��� ^9i���S
V�;�HFW؍�Ϫ�['�׀Rc�"S~��yX��o��D{�쥒�DB��8�@��xȪ�;T�#�4�׉�Y�G��i�� ]5����葝��|�d#��j��+�iˈ��PZ95����;D�R_��8�L��H����ɼ��>Z%�Nc�l�$ɐf���J���5(���dlԘH(+��N�(D��� �z�I���/����}`�}�q��ߡ��[^肠*c�z�8���ظ:�}0<*�c�|yk%�!�*�M+4f���R�z��[1蹳�ȉ�����*�,���xx\u�'�{�����
���I=�F��UDI5�j���^�)�� B{��P��P��7��G4_Y�,�⧻h�`�?�p-o1���ƟK��H�s�슖8^z�sG�`E��v��ՠ��b�,J
�ڶ�M>�%����x�������ijkk��	���J<��5\�X��ٛ�ݍ����)Ұyi"���~�o,ϑE�fs�*u��l�F]���-�F�����jgk�X��ǚ�LN�x!�7-�w��@9�
�nR��9��-1#|�OȾk��!Q�#��N2T�qz���p�åm����H�*c���u4�,ҡ��cqD�8ЍYpN�%���� j�G��e�WH4��i�Ƥbc��P/n��gD���ڣ���M�Ȇl$ӎU�Q����M��{�B���)u�2DX2��wH)�~����-YGv�k��".S��-��˹5�ӧ��n�bEy���z1/K.[����mkn�I�
�]b�M��)t��(Uр��s�{k!�Cf}�n덧�ۯ�P}lJ�%6g����'	Qi��A܇�v�ʅ��Ç�x9@�SJ{Ǉ{�Dr6���������:�kD�
Gwtxm�0�$Ex��/��ƣ#aMe}�U1��vdn6jJ���!�� ���q�a����i�n6��Ŕ>%�w`� �pE�t��2Wܪ��f��.�#�@aZðVi�O��ε!�#~�|g�P��c4H/�
��UsI��₫d���æ��f�^~iR�@�.�if�v^s��ݠ�`Q�V��� 1/�j�� Q���M�_[)��%@��i%Gڲ����C%��>�yG3ڪ���i8�M�yלv�V�7���њj�����|t���،i��
�������K��PL�Eh�K�?���ܹ;���^�ռjB���[O�J�Ƥ�K�;������8�̺7�@�[� 2s�%�&c��O3��C+�B�ՃA�V�_��3j��6��<`G3�
e��`^E����h�;Y�$��~��NAUC�>1%FR0���䂢�p��i�E�G��QR��DU���_�I�w��Uy5��n~ס~�(��nn���)@�̙i/Y��\�bZN�bc��y�E�'>o Z�������������u�%�~�/�˥�VGJNNT鐒�Í�&Atע�;��,� �%��I�����T��1�ꯗK�4�$�P����e	K��ɩ�է|/�>��q��+&5�s�:�cxTA[��ht���4�}�N:���p�0�W)u8��<�A��\��<�2e�:/��B"�N��.�<:.u��{���s*G?#��:���F'�y�I/��}hzKY�)O��@������=V���y��K����I䟨P�3�VA��ő�jf��D@B]�=������>�6Ӽv�u���渢=C�)S+����\���2B���̿!@P�x'y�WUq�����}S�ܴ��}�w���D44���Pn8ԏS���bbz`�-a�~o��(��)mz��ta�xs�pL��,���KF탺,;�����F� �ڻ�$�NP�Ll�G)A���7��WdL�����t�2��0nz�
�Hp
$m��W��}�S
�N���v�߹*� '^Z��Mj�u��ݧD��z��;��F� F�<rSE r��C�(�h��'y��Ȕt�e׷Fj6j��S|���!��&�{��O�E�S��E����},jƧz��@I����CY��g���3�m*������J[�=t �#����C��/�Zވ�Vcj8<���2�4C0FFG�
��EӔ�z4J�s�Iq҈vĬ�.���/Ēc�q}�r��'��M:�*n&C̆�/�=0�O���T�׍r�ʥ�2~���r�v�l^t˲�I0g`+:zL�}<o+��p��{�k�7���u�ٹi�V/�?܊��I���)_��)T���g����F{Tc�q�T�a)�D$��z���	D�(}q�LDsT(��ڎI���/��EN��܃@�Yz[xS���WI RN��<��ɱ����A�m.����!��G���ŝB��Ù7q�D:�v����u�]h#<�T6d�D{n�NQ�g�>LY:	�~X��a�_`반�7�s*��q �;�}�	��;,�#&�'^�Ƴy������5ķ�`�k�o�S�Ӓ1L���T�5g���.���T��n���י%�����x��ή9�:h��$]e�����7/3Xա�5<�3o_3��!{��}T�QjReu��ɳF�W~[d�������tڌ����C���۸���#��<++g� �ئ����0��O�@IN>!}�g����]�US�-+�nP0tR�j��4�D�cy��ƾوOUsp����H ���@����9��Bf"�-�{a����>T5�*�})����CͰb(�PI�nص�˷�T8����-Я%PJKu���`�?�*D�����WX6n���e62���������B�[�<\���x���+3���9ԭ	~T{)�㋤�,��j���:ò� 3��o������.����C[K[���Y��A��.�ćmA�<��g�N��=ׯ�/nn�R���ڝ1������Z
��t������)*S���'�N4�P�]c!(LY��dRLo�㍈kK�o�c9C��^}pvXЊ�9�{1�KӮ��0�$2_q�t��p��������A�_EY\�߂b��n4����g��Rf�>Jݦ�J��Wrq�rm�y����Ilg�񎺨�2H�L�`��Q������R�������]z��k�(źj���c�(ڗgq!��{�YI�X����Enr�sO�b��]���p�ψ�P���
���v2���W�{s=�$�2
7����$��	uَ4��h��.�%���(6}��p{32\$����!���c5̢��M=��O�98�ELw�2���fB��Bq�{�*k�бwF/s�s�d: �;p�w�oK2�!��x+9�[ּq�N80i�`��gݖ�F����6d�]��X�x��(;Ӕ\�5�u�IJ�v����/��! ����R�~;��������!��O5E[���V��y̎/�i���I�������|�S��W������T�ʝx#pі,7��f��t�g��v�"Vn�t���D's�ʢ�e5Ƴ�x�'��(�&fOO>Y�}�m�&&3O��C�v:��%ŕ��	��бt�,K�!D_#����s;�ÚI��cN��#<%7����mk>�|KeS��؎%�����$���CP�Z�yU�Y���¬�x/V��{�UT�e�R�T��9>�E�2������Q��JE{�AL~�#��>��)N�N�Ѷx�B#pptc)�l�5��B����g�l���Hj�#qy�/�B���?�o�ծ
k�=n2�GPӁ��ع���P�$�����A�+\Ho�A��d�ނ�g����Ϯ�\�7��Z�v�w�l%���.��U�u5Ut£ �T,�Ap������f�])!��߬��͇4<y����p�	�?�bzA���fZ_��͉�M�"����I� ��(�LF&�o{F��&���&�}-7�e���\� ���ܶ�6@�LS�r���;��'����;�N[t�Jt��;f�z8���u �������� ����ǎXm���yd{X������w�V�A0@ݏ�!6�"���,��Bˆb�w7��?NBx�X)���"��Ő$��D��1�������b�E^��I��i8�vv1ߊ��#���೾1��w��y�L��CՂ��jp"ڤ�΂�wY��W�oi����v��=Qog}0~��e"P���OKyu"2�}s}�w-�A�����O�e#��Q�CA&$�7cM��̺��Og�����o��g�5���%�e�������Y7�J����8�<U93�3x+�ʖ����ڪ��-<�wf#~��Ш�	{ǻgQᎌ�9V'�0��[Wg�|08�ݣ����G{�]�/���n�nLxNC!��Lp�^�e������p��օ�be弛-x`*(�cK�,\C%_cЩaբ5?��3�+�|2M��Ygs�. .D<8��֢�9,k�}�n�v)(�/���-'f�0}l�3����gփvDn�,6q"�	�O��4�f��vy��T%m:���CX -[[�b3X	�����o#ƻ�(_�%���*�'U���C좲M�{6��B)"{ǻv���&�x/�O��v�n� +̦QߝXC]�9 �8~�L.���A�j
[�͟]\
���R���=�u*�h�,�H�������9t�&ɭ:S�������$�q�a۟1`<a 0SѵyWS��-��ͅ���H��Ʃ�'��2�L�X,��)��i��>[$�79Ԩ�$G��q�ܚT/��J <o�"�šc���ГA"�=K�$��B�j�IDə0�F�-���(Ŀ���:~PW��Nͻy��B"���@����&��QLk����$�)0W�
�\)C�IɋkBd��Pe<��g�	��a���Qנĵ2�� �W�d���u0���i���R�&��@+����11��s$~p=�!D�[1�#r����1|�-��A6%�j����b�)�xJ�Լ��?�!�H|�D��GW@H�=��c	Gi0u�t)H4��=�a��Q��--�;���}��x!�����i0G���UK���{��i^�؀��dWg����G� 4ޏѧec����S����%�Is� ���z���!u;���x}@�=�<	)DV�+E\J�;�|]�q,���7�	i'Q�������Rr�� �Γ�E�Lys��X�x8�e��7��t+�E����R-1���t�Q��E}�`9Y��:3�,�3H��'^��cY=d��m����#@����Ј�݄��I),����=��}����v6�f$��f3�qe6y���9�1L> �z�c���6�$d�HO�o��mBk� ��h=b��(�y<W�V���w� O�4�"�-d�a!���|$�L����sO'ĩ��l�kܒ�ѩ�7��<��lP��E��Ҋ�$�TǾ>,L���FW��*����+:�a�u��5�鈔9�0Y���۾<�A�&�u*x���9��Al�4hx�G7��8�&}fJ'�2�Б���Ğ��V��<�N6���I�X�w��k5V꣘��C�0����=0���@;"��+��˭2������� �S[f.C�s���+��l�pW�\,�A��zb�k"�����Ma���'�*\S�>wa�V
Md{m�&�Ѓ���GV��5!99���!�2�H�~L�z�h�g�_����3�Y8��4�<���#��T$�'f�hfIE���z����7�Vj�0|Dp�O�����o-d��+?��h�*Ё��/.g�]x���i�VH� o���U�r�`�g���+�2cVc�TE�Sv�C��KB���~�9w柒=PǮH�C�=]E47�>{0��p���� �CA ���ɾ.�5�jP2㦦3+W�I'ZE�q�\�2C��|/�slՓ1ܛ�+�z����M9�}�?e�ѵ�/4�b��(��B� Z>~V�� �i�sGk�f.���K"�uT�w�l�5�{b�_���+�6�i�%�hTwWM��F�^�ו2���W������*Ø��T�*�ev`����t��������R�t�ի��@�b�4�J���s���ݻU�V
�A�j��Eh�~���߸ ��������7�w#	������/��٭*���+n�+$} 5�@�U�~���E��5~-�j�BM�7�����=�GN����!)�d��q�ƾ!H$�D��?���C����f�Z�^�a�ۭ�	��X�6�h�f�`�����T�n]Un��]y��y���	]8���5#��d�d��c�C�3Ĺ�h��X
O���8�~��u�+�����D�Å:yuz���pI�R�����U��jlWjI���_r�UA��ɾ��u��o)w�cf̾#�	E����|�Ջ3ͅ��*
��DmM/�R�[���	�Y}�7�%P��t��(��L�g�{%&�Yy��bt�+#'* ���6'�C�p��v��p���L�)�\l2����&��f<��$ճ�0�c����\_�?ՠ�w�e�Y �Z� Q���	XW�	|Y���s��-�����l�8 ���"k��4����~@@K8����/�S�\�(�_B��b>�M$|ȏ����Dv�=]gbZ~�{A�-�C:�Po4�f�2vt��R&��E1x5���_�o˻�p��b��є�ƔH��a�Wvq�?B�h.T��&6���E���t�l�/��i4��}���Jj}�`�t��!:�E5��j���D�Y��W�F���k�X�$}���LM8�y���?��MŪ������ D�P�ַt�`�2������ �p�?yP�՜��5�Y���H��@�LV�ٕĸb�16�Zl�^j�t�GV뱠Ŀ(+�F���3��Vb�!.�屪�Ik-��n�E���zoX�N�鸤=Tm�����D	���Fy�Sg�kuj�F춀��Z�݆8��頦�-lUZ�zbԾS�"�)�9n�hnk}7��$���9P6�3Ȭ%�v����]?���9Lu�ت��SN*KZ���#��&��%�xw/u�I�����=���Q� �l��R�(�|Ѻ�in�bՑn�duɿ7�4%e��\ˉ4�n�[�6Q��xX}h�K�w�T�fX�O�������7�v����X;��(C(�5ÿЬ2��ޕ�o��G9{��t�\\,im�t����y�z�M�蹆)k���B�d���MnT�b�S�^��qm~���M���W�pe�������O��>����(�˥�t�o���\�s�A��9��7'L��냌����F�q�aG����|�C4�dd��i�3�ǰ�4E��`�h\�;�@�a�ҕ~q�裖g�.��󮧶��Cٙ�)IasZ��t]��$g�n������ ���G�?V����O"U4>p���Wo�p-�l���1�H[��(�׆���AeE?u�DQ��"Yf�}a���Ә;����!ziL�I;�d�C8{o�=�7G��O��$QN����c	�ȇ��ܗd iAZ-��g�(:��8����,��*X���	�פ��E�������j0�-�B���Ϊ�{�<����w峸�+
�٧b�}%�V�p!��RKl.ad0���/���wI��S����X^�#�z�ݬ_ �Tf�w;KFe\�pZ߂4\��~�^!�S$�.�Uy>�RT�I�c�}&�Cʁ�o�!�L����a?9c��u����a�7+�j��Ѐ5ܣYF�`��V�nN�ҮǇ\��g:�cE?l�J��W�M@c�ྭ	���Ġ�&J�)g��l�~a�0�Q�
�
k�����B�6�u�cr�T�"䍊E)`0������;��^�*�5Y?��\���W��5��,�q�.���\�c�d�lW��}��^U&:����ٴ�@��9�M�f�0ْ���9�%8��� 9��!m)&D��#$��0��"A�RH��[�R��+Ѷ��{cA���� ަY�]�>�1�Y٤8C�>'e�5Q=�J�:��8�tS���o(R�o��R�e?6�����I��I9�N��.�߲
��n՚h�nt�x��0��Hޝ���#�04��'QW��T���MnL<K%��Q�{���8���1t�Z0�y7k���-)�?�F�U
橔�U�š�b�VQ�M��oR{��������]���FJ��&fqIڄ�z?m���K�3�^�g���)u�&��-��)�=�~�t��Si�9 �|螆�tq+��W(��/6L�1E0\��&��.4�]h�b�{��8Y6��cO�&o~/!Ε�,��a¸X�8�tƬuF�`��h�|��qz�\��A���M�͌PL��c���z��tg҄`�ծ�n���#��B����K����Wsԁ��A�#�씬m�;�wcȅ�,O�a��	��(t+?`�R���� m�"����̹ީ)��O�?���^F
Tɨ� �ϐGX��N�8�l�%�"�~���o"Pxvvl�P�tp��?�1bcx	Ǌ_p�˰��,�M蚄���(���~���w�%��3p3������Ζ;����{��NKM�ő,h�������;�4m�h5�oZ0s���דS�nƀ������LM%� �֣�y��q��GW��ڋ�Lp���r������_Xd��	�`�*Oϋ&�h�DR߱ϖ�K��:Q_���9��9�U&���6�1a�'c�������,|-��XZ����s�ײݐ�n�TAʻ�� ��l� ��t�:
s+��^��G��M��mt�R�0+����2�ń{Td�_J�=&I��Fb*ڮ,��6X�(���K���XxZ�Մ��2��,�L2N:gK�oh�-����l#0�D~.(�[�Bێ��b!zغE�i�tKOƂ���K�)M���Z���B<�!{u�ĕ=�:��Or�н�	Ԗ�ї�Ikiĝ��˫��U�L�.��l�>qC���ˢY���Z����Jԥ饑P7h,!l7(�u��R����d%�y�	�L1Rv� K�����U�4��`ev�Kk`��Y��S�D3���
-��{�Q�X�! ��#'م�,�..���\�< {3ܒFϒ'ҕ����!��# �4�E���#�c�D�y�����}��rOs����}�0��5��>1���#kbw���d��R]S.c���G #��7@$���p�]>�<��u�^�'�9�V���2��i`5N��:y�ɣ�L�1������'~9M�H���`�����+Dn����uL�<0&:?�lM��';��Y�T�V�aPk81�����qe���v�����w�5�D�C7O�q��� ���.���	��)u& G�+�h�u�h;��允)FO�QZڋ#�2i�I���/���UR�y��T`�9³��ڢh]?R��
�#gcA���a���PV�	�-d�?���Yu�|��l<��Ov��~��z��$`zA/�����K�({�8?v����^�a��g�`4�g�eQ�h�R۴�wn�K��<kh���F�bTP���P$�>�nچ��� Aq�|���bׅ����󅆝�e2�!h�%��2"�!�ƕ�	�����8�>>���{L�ha�A���|��0���P߇�lR'��������.�pU�J� ���j?U)���T����	������ӈ�v���qְ\����T�n�_��S���߫� RZ��WBy��iOu/�&��$T*R�K���#�.w��;غP�vr"l�Kd���c���CJ��^ v�
�˗�����}�dY�5І�{p��8<�3�ދ�&S�PQ7X�o�^z�
tu��f��QM5~k���+��K�Z��$
`֣|~� F�'�D9"�W��������|�u9VIP����Oq�x�M-���K�"������h�E�%&�F�Û4�X{�U�]P��VO�c/�Y7!1M|��|�Rn�T���.�U6+^���`�zvm΄K�)�Ů�06u�,�T�E��IJ/-xq�˄�N��F�ְ!�d�=�_�oޢo��^��h��U�:�\v�j��
d�vA�����Y��z�]׬�e�>>�t΢�wWۗF��7}2}�o���>(�d����9n|j����0tx�r�����U�!ےr{�t��J�����S�Ճ���jM`�0���YU2�gK� OI6'�:Vu�}05|�RǇ5.c<_�N*�a���i��]}���ܐ5��m�H;߿dvR>�i�kR}X(/�m��
,Չwھ�������3�"�!�챤	ՙ���DIo���/<����K�B'ux�P�B�~K�U^�0G�RKr5A�c�j6������5%RƠ�x�8����N4�� �Qx��V����Qž�"z*&�kܧ`b�	��}��#�K�p��ʃ��fR�R�+�P�EU-�!�`�B����ˑ�nO�S�k�'F8i��� �ưM7]d��
�N�T,����W³�a#�ycfV���s;e'.�����Dtl�p�"�'��`,;��H��ڟ���6s^�*q1�4��2MZ�^���ۛ0V�����B������lc�5|�|�~ι[�Hñ���փO���0ODT�)��0�&��T%���2u����O4u}���:�0jշ>������j�LDa�:��[��J:-��^���б�Yn M��"
O�R��g�:��le:ݜѦ4�A ���%��+�����Q6�L����u�F��Wp*'M"O�~��"��Ϭ��PCO�z���^'92v�g�P2]<�ד���M�޻�3A��Hk�Ωpk�o��p�_m'al"�@7B�:!�w0�{FT2a�iK�`ҴB?K��D��KV���@$�#�n���|miA����I��ǅ�9O:�G'�c�4u�lgDȫ��;sM��ݨ?��x��Ep�wyIz"p|O|�X+��� �2g������~�j�,������ٓs����Z=�{ߙ;S����b��گ:;z^�:i\���;�)4�9g�C�Mu��h�;��~�bv�6=?B!����Gu��lY�YM�ԨOi�39�]"c�
k��%�o㊎Oa���~�p��jh��a+��u�4���<��C-��P+��2�B�z�Vl�p���&�ki�[�l��`y?�9��==�&���ES?��>VΪO�ڔg��NƟW�^�	2B�Z@2���S��zS�(�&VO�Q�s$�}�)��'�������<�����Ũ��W�}�a��#���@9cE��Ъ��UP��/Ph�.1!�؇���V�����:DcSH��*���e9.�?����n�����^��ĳ���;3�G�5>]AT=S�]/��u��� �P|m�=�_/=,% ��Mek����?���1*v���� ��j���gn�?�z�;J�g�)�B ��Ps����`�Š�ԣ;QD���Bi�iK|
�k���e��X �5{p��w�~��L���f!� �NW�V��M1vk��οK7�8@gk#���v`��G*�]��sR��c�^f�������A�m���"L�1N6����VR���L�=]Y��#o4o��lEfi*f����J	�B�6�L����z�G���f���H	�I+V쀯�D*Sk�qW��\�(�Z������rQ��k�N��5�:Z�����Ή�y2��Q����	��lHs
]9��_޾ ����z����d.��g{� k?܅���j$N��53�R�a��¸O�Q_�8e�h���!c/>����fݡ�d^-��Ye�:%7j���&+��x�LL��˖��"�C5"L�_�k�~��+'��ΙF�c�)�N(Or#�7�3�=�]g�FN�O&���w�2C�l�j�lh,�rڠ"�͐�a��hTՖDM�=̳t�]Mnf�=��ſ�E�Z�@(��o)w����6�#��2��m2y��0��G�)n_{��e&V�n�
������B���9!�J΍����/����'�� ��zB��R�'�4���83�K�|L��Yª�u�d`X�5��X&� x�Mi$9R�U7[��R^�+ �&�~ѭ�0�K���i�4�A�U���p<�[)cr��s�t�R7`[O�K��w)��X�s�sKi�~e��8:c2����I�0�7�ŧ�����0!�ΒX3-ӍCv��"��!�f���́�R�S��bL�:���]�7��>
+�i�*1v�ɱ��f���J�ˡ��}J�a���� �^�q�=t�� �Ŧ��1�n��޿����^J�_�/�mzk|��"�^�3 �
�a�.hXl�5��� o���K�������*��>|F�N�L֔�!lA�~xEa\}n$}���@��s�)��;C���T�%��G6(��3����Sbp��w!�,��ӹ�
Ev�ˋ՛��*�AbU�|V4L/_��k\�Rۡ�����Di*s���a�h�gyW'7���T��������N<�yI��&E'N�w��ձ�%����0碾���]��C`UZVy�TȬ>�,��	���-k"}˺U��ߞM<"n��m�xL�,��f�y�h
��J�@
��t���R��b�%R	�k3��'��1�[ȂɊ�	ɤc����yM|�����:���
��R���D��fƯ�i��s.����T�e��͝�$���S���]�8CK.������U��Ǵ(h���	r�	��?���OtW3i�߹�ְ��	S�KX�~�Jq$��1�3{ӯ�o�5���h�����!��4+�a���g�T�X�v�9���)͆fm��P��_y#�|t�2��>�0�(��$L�Ť��6t�0�&�#c��e��h�,��W<V���\�<\0>:�qѽM���qu,��1!�ֳ��'N�N�kD�6c�
����H���)�̓�������~�ԓp���D�}-Q�ZϢd�K=��C/�]�AB��k����/�j'� ��������f���kf5��y�&��m�swx���08���D �w�4�֝�
�j�'f���s��Ĉ�H��8��0�{��Y���B��=�W��ʒ�eWC�j���S���R�Yĵ�%�7glv��N"�����@]���Ԙ9t?s칚���I�(���x[Q^<fۇ���8��U��|�X��Ą��<s'epi��2��G8�Ow���G7N+�Ъ:(���{��G�K��ے�3�_��z)�#W �.�@�\_�a�4�Y�VI�5�xU.2���������$������П|�$��1�i��)��:�PRE�z�'h!%"`I����֥7���)u����i{�'e���Z-��ǜb�
y[���DqR�c��;��&����i׃��o��o��A{�$v�ג�V�rʖ?���ȜH�9���I����ko�+��U�?�w���$�/�/bG�u�m��?��~��äA�(�
8�Z��f�ӿ-
���!@�[�5Tv������]�2�'�A�����$��IK޷[J�4���V�������	���n��'�a	�+�Y�Ƴ}�Q��"��*k�}A:~3�0�<:R?� ]k�K�R#Ebrr��'"j���+����*����LӃ����sW,2���Y�x8xe}�^�=2p�Q���DFs��a��S�[�E×7U�\ eB
f��מ��*��O�E��0M�ohLo2�� W��Ke��w/�^xv�77lĒZ�Eq��؉ӭ�U�t�7]��������� 8*\���, e�Zm�m^��"!��j�D�$J�U)��J�j�d5z�Dp�c&����d�vV��I�W��I/nBl��8�^T�/:ā���|��ٚE���G�"x�J���t�R�ʹ�$)�Zy#��nu2��e���ʉ2��l��Ͷ�	�d��=�P�^�(D�����Q��M�;�V5�����<�f��~�:�֐��D�y���=!�
Y�Pw~���:X���.�0�!k��PD]췲����^s�C,Q���i����ȹ� ����Gz��#��O�U�b}W٭��6�c�=�TA�ރ� �1	�URa��-��
 �+:�@}�f�&ye���v}��}�c�����R��H���ܪ:N�BI�)4J��'W�7r�	���	q@�p6�����������N�=!����:`��Đ
fU�H=;���MP�g�A?r emv�&��� )���x:o(��.?������o'�b9�"Go�W��i6Y�e��E��ґ題�X@K��CЖ!�i1��nS9�����*�/��ҡ��ˁ�ifJ�k���} _��\ �+~���ԏ ��*/���RL�Nz�Z��k�Zr�V>`�u�d�Y�ⓟ9��;�ﾢ��稆*�����G�s��K!�|朐��J�h-9��|v�xP�Q`��Tyy;��R(c1S�m��q�f�BB���`ֶ�O���A3�Tn�0�E���:�]�ۍ��0���5I�J����u���!;�y#��v�:��힗�i�8��h�J�*�3���I 8��p��,�\�t��yB�φ�zV_�ӷ���j����N�up�>X_�f�[��
�ְ�P�����z�d�>���d�,#d�.ם����Bl�l�t���D�QOD>��M��$��S�8m1��Ĩ��d&v�r�X�f�t���̍�&M��Ԋ$1���6�J8�U���Xل$ľ'��թ��-�[�C�I<M�v��ry,_=�em=���r͙h 	.j�n����Nk�s��iՑ���O8�F�#����@�B�Fp!=R@'�lm�/��&q��?����Z��N�����2=�dj7�)�J��I�Jf6m��c���<Կ��@{��$O�q��ԅ����VA]��}�hA� ��ϛe��������/͙k�,�y}�II���8��V�m�O��@[8��?�{)xN�Vѡ~A� �
��u������*2�u�"�[��ngV���Q�kge�?F$����u��,���Tڈ)�Ya�ӢU�&��M�XZ�ݞ�N9��OW�GPL��T67 �KѬd&7s97�b|l���-�K�M�<-?��\�S�Bd�jJ��J�%��"��#�t��4�Ɛ�'�F�v���=OA7��n�W�yH gƒ��p�}��=ɳ~$�x��
 ���ě�_����BB�S������,M���o�*��_�����7!Q���A�2?x�o���*|J\b�c:|�\�ޒ�*�V9g͉���{�����/�L[\h��4w�g!#�
��P3��A'��oIt���z���^Ȏҝ-��Y��_vYӡ��a=:i�7�^�C�aH9���6�n�5�^�\&� �'�뤗.Ֆ�t�?�:� G�GK��rotЙ'Kr �=�<���V�WϠ5J��C�1�m~H�5el����5~".����۱�E8� �s���������j��8ևѱ����Ӎ�<���\#kw5j�X��	��*�A}IG=8�q�$m�߿1Is��=1^[�R���Gg���m^J2D^�ox0~��y��'�08y�k�9g��v��� F��\�����3��w���P܏�^�I��Ę�SB��[	�R���PF��v��)r$�� �_��Q�:L)�M�&�6ŉ��7��܄�/�A1�%��3��S�;�UMx���%��%É;��`��'��������y�#{��;8A��<��(Xu��6�%4�l�S�VӇ�ayY�M�
r߽*� 9�B��q?D`�Gat�t�D
k�j��=�p��wf��*	��ND+n��F�tH�ѓ
D؍���(��,$�O����t�D�v�cQ8}��(��n�����%2>0���Зw��&��]5����ܖ���n�~����Ъ�Q�Z�4ɮ\�x�D[�0>Y4pTv��:4�J|T�e�6��ESF���v,�z�ȝ0f3��'��q��v� 3"�r����cf
Ovx���yB�t���&Z{]������ �=��<��~Ё��i�K4<C+v��&�<�,���CWUܕ�f#뷘���b�7B�7�&![ņ��2�s/��/9bO4U���֕�
>��Ȕ��&)�
ȕ��ڃOd�7��:�,u��V����:�\*n����t�Q���Z�zb*�"+-ʯ��]%H�����7��������J�Ϡ\���1k�ӴYͨ�*K.3vI��ɲB��vvL���R��w�-W����:t��Z�Î�DZU]�x�no���pwq��T��AV�{������L�Y���\�G���L���N*|w�<y����P�9b����d$m89u���!�Q~�6xs�HB�ݤ&it��=�ի6� 퓴)e�*��{���V��bR�S�";�j��1�UI����v�� ���$3߳�ى8eǩ��5���)<�K6ҭ4n伣�7�р4��`$�Fn[
+�n��~s[��0GG]�����8f֗�}���(�xG�u�£ߢ��Ek�|v�#����xo�ǝ�~_���*���'a* &a�0:C�$�g�F���Ȑ��@�n]�ь�]|��'u�N*\OB�I��C�#���̥-5ē�p���iؠ�v����`�kl�.�f!��J����T��h�8����f�l�kQU7�p#L��`���F�	��PQO`�/3/��Lk�}YJ� Ӻ7�&�f5�miktx�j���p�ic@��W8{7����ዯw��fU~�Q�|�5�=@i�碤"G���Ih,Ҧpu%���0�.7��=j�G����g$��ˢS;���Г���A�6&���8�,z���[�^ʞ���R1E�F��vX*����+�K�/�+�I�CN�z�kU*

����;��*#@b<�§�,s=C�c�j^a���X��ԱGJ��9֭Ӳ���t�n��MF+J�1��q������c̵�n�L��8�9z�85^q���2�]?�+:h�hXzct��4��c�w�K�a���˄�qXl6(��y@O�\�U�¬��2{Z�i4�"�^�h~���I4���ӓ{��Qn|�C�C��<^j�fmlަ��<���~�����S~/��[�l��@��2��]:��K8T�SZe>}Q?�w��IZ5��c>��[Ӹ=�]F�xS�݉3��X$ES��V���Ubb �"�H_���ۜ[����5Cj,<T��� �����w��fݗ��Bm�%b�C&Ӑ��r-�<�Pm�2�~��r��}4�ɭ�`c���M[v�%A~I��W��Eb��c���Y诡�]�bU�"$x���՟#B��<��E����F�{�s���ז@7����*5O��!-n�������ގ����~CM��(�F�,�e0¦�NI�����$2OtBSʹ��+j�sL��9�h�}�p?������ݜ��gχ����N�h�I��:>_�,2[D@�����{��m��E����3#q�nd6;$�8��+&��h��%W(,^�>}���U8�E���/�F��@̚�(��nZ����K�ش9�t��,٨��r=��F���]�����]��x�4�q8����Y���"��|�̐��:$F5;#�U�}��cώ��(%�c�
�2�.J��Vk,�N�R����|�k-���ͮ�D9K�޴���"�(���k~3��d�L��5�ٓ_��f�.<�������W3�6inZ#N��NW�Y#�eo����NR@��\���ۯf�0��>v�N��,p_��o����{���q@�7���?���$���5�����3�=|��7&y��N�p�~�q>V��=�u|����s�pL��/�1�6��E&I�>�0��n��JU��h	����r���[������zů� �̝�P�����l���qWb�&�ur�'�	���jv��267`�^�%��؆�Uh1�!Fi�ߎ��poۉ�|��$"|�W����9K�����'�[@=2^� O���X�<Z�gP��k�pf��~�4|!2Wj]���qd���wQ� Z��� ��X}�GMo�^f��/MZ
�@���yh��Z,w�=�m��~3�M<6p�HW�z�_wZٕϖ�?: ��N�R���#���oH������ L`.{(����'L��Y�fi�t� �u���D�ۜ���D}p�/��ws��saMsu8��S�Z0C8��~[hHz��\�R��މn��2�,|# 4���<m����*y�+��u�.�����1hX8�$�G����
�ц()��	kU�{���MR��ܶ��~�;�4.A�=Ǚt�7�?��,p��|�M��
0U���j�a���N$N�V��,��=����[�Xlu�g>�J`S庡E�{V����������SP�~�����%.�9�]Z4��Z���$˫�mɴ �|�k3�.��f�\��i���<��g�eq}�)�׆�˅�W�hBu�.7[�?0D0߼84���l�Gؠ�	M����,D��	��,P�v}F���aٻ��r"J�㿳nu+5�c-��WJ�?}��`f%�M�e/���T
��>�+)�jN�}����Pw�Q�2�Z��X��@�����5���K����BVw����Θ�6��C�-�iS�g�P��m�$Xfk�E!ii���e�5<���H"�{�ӦĢa�H����A�ܳ�Ny�|��j�~N���q�K�;D���5Nu]��a�z���#H3�1��`鉹�s��]�<תʺ�D�U����*��n��n�ƽ�I�1���<��A!/�x�a�<Cp)I�EJ�N_-�@�oz���9�<�E�9]Y��*������gI����_��s�.�anuԟU�]8}�7�7�2��_9J|���W����2s�px��wʮG!��;o]�a��ǅ��@�Α�C���i���_3����q�A�`T;��2g~&z���^���3�LQ��&�� �kL,�I�Ld#�_�WXAI�]�L�O�8��_��';+��k��6�t�X����ӣ��Z������0'͝����I=4�TkW=�S3ԋ�c"�1���Y%�٠n���O_�6bgt���/��`�_���U����)�z��� L�Zl_\��3�*���pTo�uLW�a]��h~��ha7Y��}ls�����ڈ�;�D��v݄@�$*,e�"��]%��,mnf����=�g�����E�gF�KR֥���K�9���j��t,�+�w夗ٜyw+f���a�a@w?X@V(�`�Z�>����k�è�<��45}����7�6 ǁi|�1�"_t=�㋻�W$���l "�cQ���r�����]6gb>�cC�k�B�8�5�B���p��`�kwZ��v�H�9���]i�������?�L���n|V&ߧ�^����M(Qt�:���F�C��h��� t��U�Cb+���������ka
���	�@�!�l��݉���I�)1������Xd}Z�Ŵ#l?��w��PY�rrT��G.d��pi<��d�F+�&�$
�cNK�E���|���2��/�o��7DО������T����M�z����daZ��h��
=��-6��%�@��
��A�+^4�[g��k�\��A�Kߛ(��'g���zM����IY�PB����2���\�r��'kr����k�ðBȜ5�{��=�/�N�BO���Wr�C�Y5�D������i��Cc�o=��P�`a��5��TE*�_��r뜫ߌCl�۪��Eo�����LaY7d��������vYQ�x8SA>Q�e@A�C����z��K�zJ�ݠ^?hG�x��b����ìy
r�;��9=`�{�.>�F�%��T����.�v��g:f3�?;!�ND�~�:xt�m��t|�'7���=�[�[' �G[R��7I�PVd��j���J�8j��j� ���$?x}B�<���d
Ŋ��� Ǆ��0"���g���C��0V/螄/3�Q|���ɜ���"��6�����]�-ߐ�d�a/��>J���M8Eb���d�i{�A���Z�K\_�X�n�o7޸�+�2Iol����ͨ�V��cK����~&��������:�R1h֛_��Uv����	ӂFz{��T=�.��W���i~g���xE�tQ�{��%lV[�q����n�	4�B'g�s*��l�����o���H��η��!�IZQ톅q!�
l�Q��V���UL�X`���:��O����k���_Ҋ��t8b<�_�^+�3�&�՗��+[��6�A�2:52��O##����	��¯X����ЋE��QB0�A]�>&&,���*ʥa�2|��ڂ�Iξu	��S�"����E��Ҩ�ݟY�xH�4�7fD5��Ө���񹼛��H�i30=L�}�O �E#�:}�-�F����f�~���5;�)��m&sL� �p��B�t���ǩ���s�MG�����*�M!���ϫ5>�"[�m����eD�I>�%Z$֡���
���[��{Es�9�,pm�Y,/�s�LD�[@� �Jՠ|�;��4�Y���i���W��������cG	��6J����h����\	D�m'�x�|\p�C�� �}����`A��ɏ���������q�t�j�L&?d���X~O���d	i�.���srϧ�c���fS�7j�g��q�d�M'�6�3�\�$���_��N���%����K-1�5���w$b��W�ݕ�g1���Va�	Ynu3���dq�z��<���Ļ�Ή� ��L��
lrNp@/-�<qq�4?���R�2����g�?��;�f�HV;S���Z�G1>�<\5�likXn��x�O���uo8j��^�S��	0|#�phY��I���[3aէ|	(�*|�����-�J
��Hl�4�K�r<ݶ6\���%���T1r�;$V�n�!f7�Ig�cK�Տ�`�WBE�^�H�q$Ƕ�0�+�B:<<f�shx���%�Ye��*x4�Y_�%�"��ڠo�;�h����fS���<�w�6ج��V���E�u��/}�� �T[�3�dj��$�E�p!��I�����96k$�n೤���O��Y�-���{�é���lQN�#݇�nƾ�����Ժv�M'�om_cHA� L�5b�Y��C3c`��k��%ã�/KW�6*��@CD�T(v�}m\�r�w�;��p|}[��%ԫ��id�v3��#L�����s�JF�%�D��燢����#��.s�\�}��(tմ^��|�d�0�o���ky������ty� �X�d�"��B=}�sp7�5m,u�P��M�G3�룟�^d�+��Ep�&~�mb�� Ѡe�4Ɉ��
C�@�n��˃�ޯ	�>Q�GN`�]����&�;m=B�G�R�;L��فI�}���ijP��B�9;Y����.tvMc#=�ʒ�\8�ǅ�E3�0�H�c̡�5VT�m�'L�)��"���4d���B�.�׭�b�E5��}I�[��`�2�C$�����Kw�)Z�T ZǿT|D̛n�.���}|��IM���I�/G������ew�N'��X���d��]?L�H��NI����'�%��붫{UߜI��K�7ӗb�����a\Cf0������:ܑ���Ww�Qw� ���
ug:�)���/�jj���Գ��>���M+�_�����Y^u�턹`�o2N�f?.���l��p�3h����Vm�:V+q*͕�~�[Kb�v��l�	�J�/�lf�m!��e�0�)Y@
�䘟ߡ
�L�&�`	h�m�#��W�C�ί����U3�<M
�+����oQ��v��
"<^�~o�hK1{Ќ�Uaj���9+/	[�'&���3��t�GŘ�TN�L�Aڰ��ity��7&�c���9f���2V7t���j�-uh0���T-P�i��u6Qr[�Ն X�Fi���q��d���{����v�VB���)��q��	���he��{�.ҏaAE�@Mo�&���"�%����e=�l��ߊ�ل��l��M9h����d-���0�����W�k�p�Ƃ�hKFJW9�z�Wg�S��% �Wu]����R<&�3qΆ�
T�X���44hӢ2�.�����W��%�w����%�=\�D���]�2�0Մ��k����ܟwKW˙kV��1XR)燐��Ѫ�N�S,�ę^��N��h�eq��c`n�H�)�k�{5���|Cuqp5��,o 9��ҥ����Z�c��i���ST�\���D.�bְ�Cm�v��oթ�B;��.ԧ��B������_�0�mp�C��MOKy$���r��ߘtS���}��#�)���U �0E�c�R�uaP�#CHv���m��;��s�����Sʜ&�*�\��sc�*�85�L�����P>ŀ�9�!�g+һ��G/�,�>7�D�"���_0 q�K������c
O��1 ���Ԯg�8�B������x� !�R8w�v�=�aK`��m\�m���p/z.�.(�Lu���Zs�!sи����_�יZ�G�P֜���y�)����B5���x�Զ���L�����,�m]������|$�Z�ݎ�wW�#��4��l�O�)P��M$g�e{�z�|�Zx�@�|�n���B��V+݅9JZ�J��=��o���!}/���Ҁ;�X Zl�6�J;������w�L�&�AW{A��T�ڋ��W3�>�P7Hv�x�t�ݮ q��4$P�O��'��v!��ʘt�u�c�.D����x&���*����Ѹ�ᖓB@���ȏؑv\�V�'A�'P�Z����S��gcd.��G��H:�=	�x�~w���mh��N��n#��ґCm�����Q[�mt]�v¨���1Y�|G{�,}	;�W^5���b�i�g�`����ho���e��V�\o$g��R�~�nNY�CD��AŦ�F]�}��ik�j�_c�(�!��z�H�u���&W�ӃtТ��>�Dl&�ux!6�Qd���WĒ�|ZQ��2vEQ|�x����u��4^�T[��#m�*�{yM��NT$�o�ɴ)n���.��͛�z͓��1��>�\Ty�l;��18~j3=m�W�9u��f�ח=���tr��
2�)M�jU��tbB�~,6�{u;�2@�:�d@�rn��j����M�B�>�SU7e�ci:��z�h �9����\���E|�cϘ!�T+2Za�?nN�B������*"���o9Ms�����`��G��֩��)#�_|�s�ՑG{b��qH�GBp�0���p;,18�'�"����m��ai���d�f��bzP���p>m�)���Н��S����.ډU�YFA�
Y���&�,/�꾹r\�Q�5�������֘�A�|)�[\TV�ugg��
����o.<,��C� ��oMi���B�́�r�v��<�XY����R����U��`�y��"UE^��lij��-��KŶ�����|�DI�b���)[y����,�,Pz���U�M\s��|WD1&_�I>��Bi���"f�~�6>!��i�"2�r}J5�ڄv5Ů=3�nYPT�g���W7�(^���.5��V���˂&$j {࿱�1�v{���(��]7vB���#J���+�r�5��<��w��u�V!��Q�L���"c
c�}�C?��Ks�n�ڕ?r��jS�U����J+�%XyB�v��8y��&��w?���LP�3�����0u���z�f����fzN�)�8����,�U�����h�$��8`i6�1��\r�a|_�S4a�,&�����z?���
l6X��C�9;{[��������Zf ���+� [��� ,���׷KZ�"
�`u!�Z�Ӕ[D�Ovg#̋�� %ѳׄ��D�Q�9����b��� o�EǙh��Y���&�9 7L�`7L�0x�m1v<�%{\�� P ,�!bD�u���o����h8� w��Mn�� k��'}GT�Qm�:X��%���d��7��"c��Z��>���ӎ��^��k��p "��AV��!u�8��^!pG��+����X�~P�����Ŀ�(m&T2z��톹B��9a��;�u�^[`g�m�����\[��f����0��������&٣/����x@D�M����R��^ȷ�ݽe���Mw���胸op,,�{�O![}�k���t�D'�|x����P�v�y������Y���I�Em
33�6��F��0 J��\�b���./�'�܍�W���%�O�O� �.�Yb|�Y�l�%q���KNSfa�"��iL��h��摆��O
B���χ*IZM��3c?}ghC�h`1�e�Wü�|��f03y��IT�&�6\��ZSE�?�:��?����DDS��WS�.�R<�x�̩?���b\��p{���!Qk��㞛��g�������Wύ8@�⽇/�$Sl:+3K��O'����|<���k�|��l�Zg�I�m
e���KM�AM��$�ⳔF�4���6\�"Y{lNl ��G�	ٯ�����V������cU��@V1�Et�z��%+U�iU�K^^������AG�_��p+=^��Q�:z��8��ZnOS�bG8��ZC#!����{%�u�p �/a�N�*s�����B�ԙ>���j�r�<�n��a�*+?,!�*���96^�G}@�����Mt\Lp��h5�ī�0�����Az���V����m�}���v��DL�c���K��ذ��|S���g�:щ���L��ռ�����S�o�HG�H������_Y[J���*0p� :`�:C2��E3��T�EF��V7W<��r&��1�erv�%Q�䲝�~��X)�įfm*��,��I% �n��Z.8./I�qHfW���c9.�U8m��3�8ew�%�㺔R�Д���Pܓ��(4	Ư�b�t�t�u���3lf���k�f��j;8��Ȼ3�A��|`,U��Anpa!{x_�O�rJ�[��W�8�s��(;a��΄՘���a���f�WWV��bQ�Jg�e`C�i���&)��ӰV����%����X��Uj`���u�����_��m��1gVyȼ;盔<�����/$H2��y%������Q[�}��[�h�L�m�1�r}+Auo,ȷ��]�o ���[0����T��K'����A��T��o�8�/�����B�����������6�ߑ��.�+r1ў*�SK[���2s�ґ����6�a���G��|�a�u�JW�ҍL�&QM�/;	¡��.;�{�9�sIA��h�	���B���yWU.��:�j�T���L���WTX�3`a�R���M�'��U���|c.3H�$gFՔ��D�գŒ9O�ˆrgk<� ����B��W����͋g( �����Y��\Cn/���DA����gl��Ml11�|6 �=��g��m��`�Z7s�ސ{���pl浇�KŔ���F��w
�[T$��v](giaM����-_��k��Q�ѽp�B=�Ÿ��z0�ŉ�`�7ov���!���5�)��&�J㸨\6�?�j%i�f�^ڢ�$���MƗ�*�!�?LeB4�;h>X��ѕ$
��#�Ħ�P=e�L�?� Y$����O�	`y�x+�E搑�tO�&P�IHPt�>t�ʄ荀�q
�_��w��М�D�=]�Jv�j𕳩\P�ʕ���x7Q՚��D�| g������h���������7 ;[<�yB���Ep#>Q�?�}��J&�!�tb�
��4����u��sB�U�QN�!�ǀ���芈Ȁ�T� #��L��B~p���@�f�7H�<Z̉u$N�R43�����dR�,��mrC���������D��̡@�B]��-ό�S�)Ry"�{ a�i�dfp*kt2@��[���<�9�[�9UqQ:H�J1;��-�d8���j=#Mn��)�P%��)=�����˫�k�|�y�r���sm�GXu��<J�'oΚ*Ŷ��ܦ�z���c��v�qu�/�"�$V#BVFD(��7֘~�EI]{H��/��4��R������:6o�m�YYt��X��RO5�l��_�$�-��A?���yn�:$�ˆ����P)Dy����!��WJ<,-��`I��F��.��ĕ�Jy!:�G�w\9;��3�ޑ�l�ۉ��P��e����;�ql�o��D��p���cz�Ƽ�-�R�2��<�~�5�r-o�u�^����=AN�"C�Ì�XƑ�Q�{|���K����SyR�a��H��[di�]�;$%7L9B��u>�;N��?4v�Jk3��5�Mf��1�;\x}�z�2��BUju\Z9'�#�q�<�F��ti�I�����ɹ���v2B��	����Y'��Dr*�0D�������R\m����!�ؖ�wγ	N��Q!sM��Q��:@��
>yW]�L�(��O�	x�xD����$�Q5v��/�@���F�"�4���I"AX��|�(+�	��g6w�^�{�a�f�l��[�d�Ͻ�9���O8��w�?�E�H|�Y�{�^�̶�
�����\���o�5���*Oy�a~J���nN�>���Lz��H�.�;+u1e��iy)M��Q�����[4���cl�]o-^�̝�!C◼t�=&�D���D~���H�z��vD>�g(��4�x��,`up��-��jɲ�3Y���J��:�D᡽��P�\Π�i�z*���u=/ʾ3��^Rv
�4�o(��]�[�Y9˹�F�GT��GXD�Ӽ��t�0K\��Y��4cxQ�Mò�e `���DD�+�W�z��b��ڞ���B"@�N����G�Q�8&������ZPI!T�R/4�J�i~�[6�l%��?������P^(DN�+d��$�}��q������s�:�٪�2���X���Tt�0�"!�P��������D����ưB�v��u���ki��MԮ�ȲyH�a����J��?EJj4�"�ġ�gA^���*k����Ga�9���n��@�(��0ˆ�K��f��,�F�+Wp����c���DBu/d��
3�k��+����KD�t��Y@F�+���pߒ�0���耇1����q��l�o���&9Ӻ��(`�ѥ�K4�L�<�zS�x���&�7*)H���U���!gX\$Ř�R|D��S�k<�������c���{ك�!��lt���5�Z'������P�(_�)�[���Ψl1p����W�������Vh����E��b�:N�=V�=ui��vk*���"N�����Ȳ)ݐ�$��V���+w���!D�e
z�g�Q��{3�������?�g#��ʎ*ӥ�A����!o@�R:\�����8N%}�n�X%p�J�st�I�"�	O%QZ��I!�_�X�jV/�'���B(8l��v��0c41�U���W�[��奖sv��Eb�i+�9�Ho�T�s����{��L/���#Sz�a���2	�(�ݗ����/����j��)�k;%LB��9��D���5�e�KAr�(	 d�&M��d`I;�|�!���o�CP����,�g{��C���g�c�ȓ��%30>|K���������*e�Dx5
Ej���Fգ����E�����A������K��Q_@b�%���\H��O�gjv��)c�� �F����=�����;��jP�����%���/1Ԋ���C������m��!�*<�ۇJs2V�8�3��,_��P�pN���7���*j�X�q��1m���Z����H�,L��Pu}((�#x ���<����+/�|��d�[�%=C2ȱ�R��M���.Kڽ����N���1�b�{E{��$<Ӧ��e.�4��'3�y��k�f��xY��w��o�=��*���y��?)׸Xa32��ׁi�ׄ���=�,���DA�Ҽ���rf �w`=y�3��UM��z3x��&U)�%O��o�Q�12 4dÿ�Q�(*�-�BVx����<�Y�V���_Ŕ��e��4���D�d� ���G.������h�		�x�QQ?���0�ŭCн��X�&��%ً�2<��}5״LAo^�N!�í��*)6��dV��R�_���x�j�2�F֯����T���䅓EQC�|���*Ҩ��)/��v�ߐ��D����R7�����}q��z�����q�`|�V�<<v[3&I
b���^"P?��`^Q`	�Tq̨׉�mDWu?��%�9�'�KyQQ���-F	��.�A�Jt,ƋW���N������7vF�%�}�����8�ݮ�G�e�;�:���[�K��iM6����w�EYhX',�4MjJ|�ܳ��� uߝEi����u�є�W�>��ׯ{��g���Q'�a|D�����&
�kJ��l5!���PF�G-)�h{(��tN}��C-#C|��9�x�TS'C���	��6�Q���f�M��J�K_�B�L�s���ϐ���blHX �J���7��t~:8#Ԑ�����.�u�a���DLu'�Ƌ^U$%�u@!�xG<��ɳrVz��� E!��?ؚ��['p>�/�N�|W�^X��vτ<K0�Ap}�^����a5T�D^x�V�����Lr���ufE���ٷ�.<a���%�6l.�7��\��b:��NA������)��EӮ�Dg�&i��U�e��1KhvAQ�e�U�'xuL�,8������1�i�6��*�/�B�Tx��M��P.<-�Иͱ2�\��=#L3:�Ǽ���y�C��	�Tb|�M,H�ܾn WDFb�su<�OV�k�:��2dĵ6M��r0��*��l�jf�n"Bǰ٘��0J��y��Κ�N��_U�0�=������b/�9E/��}o���a���֜����VO�}�$ɰ#�ˣi��MO'To@i�� ����Y���MI�q������H���vBB������[xFx��3%vD���a6قf(
���������Խ�MM�Β0�E�'��vM�-լOZ�5ub�Lv��v���K
�_��7ATQM���V�!mM��6�{��`\�`�L��O����6��,y���5��z� y��������w/(�{D�y�X�w����>�R���B�E��;p ��>�r)b�w3�>Z��
U>�r�5�Ͼ�N@J�\XʙW���i0��~��kI�x�e#xf<ɱe��VV#��m�C�L��ö�FL�d�A��-,�p��b�U���k�K�ka�EFT����
AǇ�ٕ�#
*�����׏�H��$�����������tȄIgv�9�-�U���I��/�.Y�t��*E��i�rv�[�QR�CK�y�"{�]����ӿfP��'5`hUA�L��9����@�w��sO_C���!���}��A����hL�E|�rf��.�0M���q�dAՎӞrGv9�.;&'rp.��y{�'ΨZ|5 Q�?0ե�}�=�,�98>�����N��63>7g�NN��]� ���.=�?
*?P_oךD�^`#Ys8ƛ1����+�Ȏ�j����ts|G��h����CN�S��󇂘�<U���v��2�]� �g=�B�n=U=���J���7����)���m"�T2�������&xr�w@.��TC*�� ���2���O/��Ab��� A���
q��(���:�Aʤ%�'�����u	��O�u�������w���'<Spon�#wx����(kO�e�POi1��N=���{]�Y���Tl���*$��:�QK Kpy��3Gj�Q]�I`qVg��(��hT���X����A�����H3�k?�M�1�E��h���^��t`B���f� �_?�>C�mQ�������.P��堌��|�n�����/W0��n�5�y�
HJ�A>՞���f=#�P���g�V�$`������4�n<�t������`��Q�v}jB�gd���E�e<$7O�a��3������8�ݭ�2�U4������r�� }T�B��i�%�F���x�s���F�쨙)EQ��=�߱�G\���W�� �\N*0�aE-��P�<�4����MP���c�L���A�!b=�t$S��b-Ƅ�/C�ns�ۓ�/�����.  �`}��߃�o���-����_�TA���������^�H�d�fx�vX�Lݳ��0dFWT�a���J�l�ɻ�������0��Ur��c'4�Ӿ��c��1�q�-��0���\�\�D^*�a�cOO��I�"eGO
-��_�`���N��tE�0����������Ai0����8��Hա���<�C e\ָ��ߍ���=9D��Mg}�.I/d����h�M���8\���5�kH��e���B'��I�9�����s0f]�X�d�C3��c*'dg�q��=�K�h���ms�Ιf�_������"��R�$��P���K�l���f����B2Y����V �r�2�po�o�,�rI��Zz�͖��3��׈��փ�������_Q'���5 >&h�2i��,i�?���!��_%�I]�����s�ҮiTX�����~��[g��<��l#��8.=G%y(3���2�:�j��aď��������G�&���[2�R�;��~5N��)aL�_��G�6��X k1�E�V�á�5��s�X���q	5V�V>�N�NvR�� ��Q��fc[�q�|7��=7�������VɂͤV&��#ӈ�فT�H�x�P�	��N0QM���۽���-�OE�k�Ǭ�
8!���ɲX�����`�l������W���j�XW���◳�j����	�u�d�	g�&K���R�{쾽-� ��M���œ�W*��[ΝB����$a���{L�hq������/O%v�'Z�� �����6е���>n^R����C��O�&8pZ�,��ֳC�e�`%��)>����\`t�eJ����'��@���ŋ���i
���u!�zg~�eG�]O���m��U���u���e�lR#d�o-dJ��Sf!_�6�����?�O4o�t!0aj?�|�d�Y�<q�z��pR�#�A�f�8�0!#1W�ŝWQ�F	��Z�9AQ
�)��/8B7� }����<��\b��zi@f
��1���\���G˚|*ꉃ��$�Xh���e��
�'���uI}�/ܪ\��/<�Uh3� �(���C�U�aR�l֍Q{�w��0hF�Z�M��퀨QToݐ����8AG�
�1z��:��k]�56���b[X���j��@����M�i��ҁ��^l�z�g�)>��op��zl�w�P'qE8�'����tJ��:e�/|� ��։��Ĳ;_���]ߨ�����y[^5��aN�ifO�SO�|��,P��X�7�)�����teF�؀@K���N�=uEF��kB��J���J<_��6{��lKt�)��Ș�?�)��¨$��N�k�h-�辰y�=iG��\�n$�ٷAH��GvB\�:��b֨�~��u�Aj��!�R����B6��oT����`P�������T�V���]=CR�����b��8xs�O�2L�c:���5�˵���R�"�gB��i�.��6૟����3���j�Ԫ�]!⦟Ⓞ��1C�.)�c>~S9�bg��#�����ڗ��y��X@)�HI0��.3��3�����s�G�H1\Yn�hv�ҊDr�� �\N�7�<�4 	��Z��Ѫ�8>`��[oqh���3@:�I�塇»AΛ[�df�uQl���t�2 �9�q\*]J���2�Q�̞F��Ț[�֮�ݟ�C;������LvEd�����c>��%ʂ?U�i����+��s,\�3P?���U��^�7�QUV�)<��ë�����横y���n>ؽ?$d����=���%Pt֠cC�����ߘ�1���v��o_;�<����q����#H-] �i�jU{D�����6�*��]=�+JwbD\B�X2�:�Hoֵg��@f���61>���h}��6
��H@w���J(cP�o��KU�EO�}b�j�z<fA�c���c���¬HFs�N�7��� p�L�R:Ks�35FǴ�Pk����WV��M��z�~0�ʓf@�;�k�����䲇�BB�Κ�/�Ҕ�z4\y��.K)�r�����
kq�$ �ק�?�!f{��q3�>� @��Z�x�������6.���2�j��=�`c�����7 ��n@A\��!�A�g.E\�x����-�=�����߲��U3����b$D���𾺨MB�:��\ѵ��2hhl4�,��ɯ��9ʻ���iT�ƖP�����u-ӷ��e������l�j?�x�?J��!��_��y�ɧL���$�j��]��T׷ZO����Q���ަ��C�$�?�2�\e�Y�-���}��`�X�LAV�Q�Z�����֎?>����rxIO��j�K�������@�ye�nퟀ��v�w��t�_G"/��>9ԗX��߸P��7_P�M�'�H8zR��1E,��a�����k�+���A�S	H�t��I��8]yX܉q���6�G���Y�^�v�y���΂�?��c�:m��E��=�����*bc~Vj(�2��ق^݆�GC�Z�N��H@�CFM5��{�uF�0�V�͈��p��w��a�G��D�n�J	�叵�;�A���fw��a
����(���� ��Q��2�����~"jr<�Vf,K�J���|��
�k>��������N��!�f*�4��<�T� I��˷<R �KL�'CsEv���I�0�����x���������T���}$O�d~�Cݗ���u��3)��K�+3<��|r۩0����)u˥�k�o�d���+Rz'�S$W[��Mv�n�w��Z��1�/da�(zq;F�����W4��jh:�_��V�@?g�KI��)ufQ���|
NoW����AhP��êU+�m��p�8;�_�Bg>��6�����̉�p��K���wj��V��c���5�q�X@�//'�64.�E)+3�!؟���rd�+��!�tT��������t���N_I\p��?A�>���A�.ב�4`er�\
��g`�X�}ǥ�+�Bn��3_hcXK�<aZP�!����)���)�7/2�˘������?j�vRP_	�G8���;�f"v�?�n?�Ǽ���2«�����wgo���/��e#.��w�����ٮ�:��W�5�2f��hr	�\ �_�]L���*�.rW5�ʑ�FP%�?�~:�1R$�������p�f�x(*Y�t�����D}��3�����1��<�i�,��<(�Q���I���\�3��p1��������:޹a$;�:>���30�*(��Y��=5}j�f��-�Gq���w��-r\]�iv�b���� 
����$���)���^����]1�j8��䝈7�4�%�!��J�|ȃ�T�ɜ�ua˛Q,,;��_�˥���G���9��h�ㇶ�
ώbtc%ڹ2&]�{��r��	�$s�͊�VJ��}�7"��(���c��a�P�D�?y��$D���+3K5ǁ�����C�in�1mY���}�17��a+���Y^-[-���/����_c�޷`�."D�'��9$d������4qSZSH���Z��~�$4/F��t��CeZfTz�J+�02a;잋�:\J(-ԔL
:�Dy���<ūV�����+y�<m|m�M�����5�DJ�(%Ec��SWe�!Ĭ{ 	��V��2/�/�ku����y� !���\����w���N:��(3(wD�Q���{���d�Ib\x*ﻑ*�\)T:tB�������6�i|�p��
��8�(�VL����Qe�T�X�>7�M<K~�W���V1T�(�,�%1����ǝ�^�P��7��]�j���ﶿ�;��9��X���UĽ	�_*s }D�HR�y��'U���A�)��
�wI�_�j��5π�Ж�
"�0���f��-J4����������z����z�9��u���m�Aɛ�N�l�������$�r̚�*����.C���m4v���	�{�Q!���q�LY�@$�4�ƂJ{��X�Qfؽ��O�I!���B��D>�ű����8���%��2�'��؋1��q��˞3��I�@�����܏��=���G����[��p 
S��'������f�~�������f �ܗ1<�Ԋ�����d3ԧ�-fqoԢ��_g�^|���-�q��������^!�[ޏ��鐿++��"|����g����+GI�����S�#g�^̵�wtY�h��\w�z[��ƌ�mo.�m(K����˂��ϞT.��~X��54�Ui�#u�0��T�=a<o,���)?{Am�0(�Z��ķJ�i��B�_�/�Z�%`��맔�`+#(Fs�G�b��MA&�Znw����� ���mu!_)[�I�cӧ�,���֠0����6#Qs�$=�x����S��v�PS���3B��r�v���s�8�5��v��S5�i�M~�ȓ�;;ɥXb�Yh��5dO�|�s�,�+�f�!y��\�����u��u�X�![{��b���EyC/� �,���Z���m�����F	��� ��9r�m�X5N�~����Z�<��M*7~y������M[�2F�i�+��r<�����s�l�S-x�ݩ��(_>�h� دg�{b���q�C[�2�ʮ�H����X�$m�{W�]�\u2,Q`g�JN�n�i���=�y+���P�q���
c�V��_�`��#HwWkB߮FǙ�����θU�oȭ꘾1Y�*�,�H�j�������{^e�r ԏ0w�E��EǑ�Wm����(`�w�;SUm�l%u0����&%��$Ɍ�d��T`��C�7�����T�G§ۆ��_�W0�T�[:&����Jv�W쿳�#=�����*�K�<-����^u�� �t(H����rg�ؒw��(�2���������.',��'L]��*���b��e�m��ܾ�2��Xi��F���E
@)���D(��1��{�eyE.Ш��Oo^�J�䯵�O�?�SyӨ&����d��(�Fx=����f���r���2̤�:g=�¸�{����(��t�v��f�L:|y�g�G]��Hh�vUZ�WK��0�Eo��ѯ��g�J����C}um��?2�Ѣh�~���/az�m-s�NF��aI��]��a�ئ_�;S�Iͥ�����䡇�{7p�hS�n��V�N�}�=Yv+�3	���D�N��e��l��=���Ñ�X�6���������(?��>�"Y��86(����c`%� ��b ӺR�-��X`S�*��/�Y��?�u�9b�1x�l�����g��g����+�y�!o<*���D�0E����}�_����Xň���M�x��6K�c.�{�i=��b0s�S�ɞ�NJ;k.kX������H;���&����w`b-�^�>В��Idh;��_��H��ADx,ѻ"�D��`ϳ�pdc>��!'�N�[��ek��r(�B�jj��-sN[�d������j�%>�k[z�ş��1�@�x�T(�PH�O,����u8uIʁB�kO��7���,�Q��K�w6gXR����Fp䵩���Mho]���pEs�U��d<�<�;'���4��o�&�V�ߒ��C��嗞N���U�������f�$���d(�r9�}���U���q���ȮZ�n�׬���zva _��z�t��_m�%\��P*�q���ڤ���b��~�י�?{PqÜ�3�YG��Ƒ p8g<1k8<�(��o�/-̓��#�]��&��e�������eU��XZ�bY�Æ�Eg��q/� }ʇQR.�b�-,K�(��Xd�̶�?�HoG�L߮�6G�lѩ�����Q��J�]��̊��G�N��iԠe�{��&Oɉ-�W޵Uke�8{Z��	#�L�&#��ُ���l�W�7��Kw�lT,�L��wo�MWc��w����+#9p��3Ԍ����gZ���a�����8X�W<�3�UT�bZ� �1HGW>�>���u�v/U��K
<s�"�����U}���5�[��2�g!�;�;��8�U�\P��gg��
/u;7��Ho�pD^ꐅ!�U�Ff��l�PzB��'��dL�|��7��$t���2��x:���Qb�k�\֝�}���ZWa�{�|x�f<>̄�hԴ2@�J���t�C��)�UU#�f��˜��r�G��34)�<��w�|@J�?�ܪ0��iYQ��X+GWu�9���m��tA;���Y�u�C�R���e�L�$tq�r�7��d��i\Ĥp�rU��;~����W7\m�G*bũG7�QRf�=��O,bj)�N�]j�E��n�)ğ-�G��
a�]ԙ�T���tǝ赵t�3�c���'%��� S*Dj�M����?���ec����S�8�UGir*���cj ��Z�dͰ�񙚉��\p���[XWߤT�}�j^�H��ū���;�h��ĻЃ��{r>�b(lD��1��pnrMz�n�j��f�$��#C�ֈy�04MZMv�O6�� ���Ì�?��s��ΥB�y�;�AS�-�� L� 5�^<#"nR�ȋ"���bC�-K�:�\�-���)�J<�C��.)���zv�4H�2��r���8mG*CJ���)�̫`�W�\qah���&�͛�8A��N,��j�-���
�	�x�Y���|��(�Z��O�r��莾��8��o��AT��:�r5�}���H�"���,4������4K�z��R'�*ez\LU�`���`7�����g��ew@�t���X��1N�+�]�~�?8?SF�
Y'S�=
���@HŘQ��ò�uȨ������T.�W2sQ_w1{v|<H����a�RA!Q|	�R�El�����Y�[��"7)s��P ��֝6䅦/��W�UW�*W�,��|��͉G���������v�����,!�N�������8=�����W�r5�U�T�%���Jy�sp�П���E��f�,>8�(�+�.���?�f���}��v:��W�/X��x<	�|ȹ_yv�&B�c�5'ۓ,5'��kx��y�q�����j���O�� 	iH�K�ؘ����;����$��!���x�x�=��rMv��*�:���Y��x)����x�-���Q��ӛt'���9��J�	�wbQ!����b�f��y�5�aF!0���>�}ʣ5��~���`�"6��:��gm5v��Ƕ�Bދ�.lp:��z��������S�0 M
x�S�frl�N�Ӣ0�������7��?��z�]��m=Ro}T{���@noI��� ��|�)?�i340�G�~
�g�����T͋<����.x������N�8jM�4#쥨}�]#81��x��ϡI��*\��*�ku�;��J��76xDCф]̵>34,"����K��%�����H:b���;���V>zǘ���()fL��{/8@����̻��=̳�:|� ���x�#z���H��^�`�1��� �&{�'
H�����m�K�&�Z	Bu76e6~�^F�J�HN�v�J������f``�4�ڣ�����
&L�r�v��!���r�����_w�y+�g�GY얂8W���A����|q���8Ӓu�܂�Y�����: ��k!On<���#~6n���
(=��w`?s8q�6�X����ى��N�ѻ�r�]B����yr�ʝ߮�Z؞�ك�vv���@2/:�BP�����*t`�/C�1�[I�E��4�M�̹Jn���6~��׬D���O��([���!S�|��
3R�_w��On<;�F��]=��TF>Jy���r�x��6G�uI��E�5w��$ �v�7�^h@��]2���%����:���X�^��k�{��)��4a$E!q�a�j;�����7~��\B��,�V5�>�5,�Q>E�KJ�0y:��>O�� :D�x6A�Ih�gЙ���m�m��gd�;AE8=9��{I�lw[e-T����).	�޸�$��H�׈Y����j�D�L����,;��;����<S0�_�F#}��TZ�lJS�%H7T�?�'�Y9����Mr w>�T�#aU�Ѡ�����B�}�O��7ҿgت�1��폹 ̃Rf�Z�?��n+���A��?� ��s#����Vx�Y'ac�eR5*����
riB�&Ƿ�:�a����n�/0���K�ۇ�w����u0ay�I�k��h�b@9��1��ۥ{O�ɉ���=�����C����"r^�O�E*���f���GL��q��B�G�)ߓ�
#o�
{bK�5�>0D�9]<KW�CF��8� �V�j=M��̑pF_��C�����y�Al2Ӊ���KU@
b���M���rc=�6�[�`ғ4&���6S�!BĈ�.q�(���$���9�5b�C�[:�=�����/��9�xu�4�ߑ��t���׸��J��P�sdJA�ƶ��A:��"#���Ϛ�VǢC�_��l�C�&����)�i���"w��H0��~��
���W:��i���	#qW$smS�ZH�W_V���;��R[w6����&1G���:�(F�p�I���I_b7-�c�Y;�j8��B��z6�{g���x!��u#��l8{N���(�u^\[n��π�"y�_Yu�)1E�-�� �j'qDl�;�qO�8ӎZ�]����9[1s�vڼ�s?+����E�g�&�ۭ}u^V�t���oN��k,Fx&Y�g>�,����r�Y�K�F�z,��`�iP���-0�o/W�K-��|��~ȍ��gL�R��\BF�~��m��"�#;����=��#���֒���,u��kce�D�ƀ2�ߓ[R�e����"N����%�0���;��L���<0�[�-���!F��|�S�5Q��2R��6��<S:gl<��8��x�<B���)*�����pe�2'����09���k��Rrr�;��L�s�Q�5ә:��t��͍5BϪr�����3Z+GLS��F�
J@�%ٕ%��{ϵ������'���6Fʯ�c,�(=�"��M�Ssk1r����j�{wnc���dW�����<{'9U��KF��|`�m�
���iע��"�����^e�U��E\絓/=<�ؓ!�i&b��%{�פ�~�H�k��nJ�}{�?P���<�D���w;ٮ�U����'��!�EP��S� .W9���x1b��^�[�|bڞ ��1�q����1�
��p�����A�����(���8΄ő`�k����>�M|��8�%tB�ڱ�v, ���lt曎����!b	�Z��HԀ����Z��v��u7���d J8���޸��ʭ&tu��*�E�e@ƺ��T}���χ�x���G�dn��`:�Wro��� ŧ��CP��!����>�Rҳ�;O���)5��!�O*���ID�O�h��l�)5�s4H�N[v���kHцCV�VvH�̬��X5kЪ���L93��2]��Y�D>s�L��7(N͡.;[�_�E�2�
�=Z'za��Q~������ ��&zݬ�N���� ����6�:�o��ڀD>���L���b�i	�6�#��m�։��4S�L��k���ڨr�� H�7���p�Xc�2��v�ƜuOj'�u(������w�E ���Qu��"���kYju����"@;��*�dGH�Fz�L�/��&h��>3ʗ����i\�Nsad@`l�����Ϣ2��9�R�\\����WΪZH�a@\r]��"���'�US��s�F(�ݪ�TPP
�g�ꈸR'U�xU�O��L%xLb��Ҕ7���:v�NA��q��2f�vɽ{U?W(��T��5J�~�z�qede�J�����S����*�����iP�C�5��ad*�\��[p٬;���l��íU�����?7Cr�R�1x�?!]=[KB��g���:�i>iT�q_v�L~l�a;u���E�����U��-'����?�� m����Fն�g�)�Z�;)�|����M�Ş#���j��Y��\m����5�e�qG��r>?S����{�$�bN�p�ơws���׬�a�]�`�&�C��;sC�ʱ���� ��ǿ{�K���֯����2OQ�_��*k��A��M;B^�)oJW�x��wnZe���O�	V�#�4��Z�)�̯X����\�� ��|+��I#_��s�W_`hm& q  �D���y�[w����� �5Fdx��%�_�Mr��C��M,훣n���-�z!�hã�0��y��)^��L_� �l��1�y{�<O��d錛^���0l�M=J[k[�<}�H&��XKw�}7Mv�LRXq�vDѼ�����!?k�zH�3Hm���=#Bv��0b�M�8���P�g1�����N�=x�>
Z�Mms��:�sPm�x�
uHi,�,��yx`2ͷn\{�5���~k$��^�i��-�s�+���e7�`�D��s��?dcn�^�Xׁ�S��x��NO��eV4nF�aə(�%q�����o2����<����*��?������#�d��4�U��l�M�OP�����"��RƝ��2����z����A��v�_�XT�\Nw�m�#N��8��x��-�=񟉅m%�o�V7���v= �� � j�a�	\a��� +�pc���f����	6�0ȯ�Fy��&�m���BI�t�>d��m�jw�e3H��	�8Q�ƕq�!�!�n���q����]-~��+�|�4�a�ԣ��Ig�+�M�IU)���#�#$��.mb掻�|K���$nI'�ק{)��%��A[����`�����Z� �?fe�M�]�}�}���AHGO�ہ/M-��]�WD�}��k��
���Q��7�/�
�P^B���� M叽0L��2�x��l�x(Alz՞gJ�C@��pqҗ�n�,6�ܫ����gh��~Z��o	�ӈ*�k�w�t�Go��ܵT,W	cCU8k����Jt()]�1%��lə��P��f0(h����b�Pv�F$�����Xv�m��Ҷr��Z���Њ�r�l׮B&���f~���#zZ���H�h'�}9:qܡr����?���o��$��~���Q�h_���SZ�K�@|����c��	eEf$�<C�}��N�;� {#�BZqf�n�eԚY�9��g���>���:�h`�y���Kԗ����!��ص0��(�8�ʗY���j��}zk]se�G�$h�#�O�g(�J��c�����Z�(�U��R���l�CS������e�<d#ߎ����P�
ˀ26l?�E0Sn��_�4�
M�)�k80���ve�'��͠mmF��$�N]X#
�7-����O����:Z�D���^I��}�g6�G���EEm�I�N�c�DA:��'���3�3|<���;�ƁO2q0�Z���LJ*م����j�wy�X$�ҝ*���60����~�_%B�[\��IR�_� N(���M���-e�|i��~s�#JAR\�]4�K�Q�*���H3bs���i0I��V�4�,O�sZ���Glz:U�� }WՐcM^(RO��uK��C���epz���ۋ B�ʥ`�4�1?3�an�D!��r�
�N�O�� ]��X�#�  =69Í�@B������u����k�~.�{&�q7�X^�F�Ŧ���eB�ح" ���X[���4D(��w����,3�jغ�#���o?*"���gz�*���^ߑ��d���@�Z�ŪOmo�$4W���1�kT]��b�|�ߜ"(�$�i	K�^�[}�:�Y �<�����LZ_	PT�x�m��'�"�NJ��^Bӎ�"�!��@ ���&@T:��Ӓ���=f,�5������렷o`��N�s~��W��F�C��� �ԸK����Ϥ]���0���y�4|Fg��P�9�y+m/�g�""���ֆGx+�����c뇖#T>+��ͺ����Cl#�����w��w�V��B
�ʹ�ͮF���4f$�%ژ�1G�ooG?S���h�j[%,_�F��)9|��M��O�=u�����c�K��A��g��+���[��Q����w��x� �\�
��aa��B�Ю8��>�e�pؑ͟��)��X^shE�<-�J��C��J����Lmo���'�� �oc@f��L���~��`Dz#Y�I^3w*?e�lPTY�38qU���W�5��+ �ƶ�\@�O��w�|�⌮s���{�%JV�T!wL�'�X	9KYJ{�aD�:�v8<Y��j����Q����b�������V�Ī����Cؿ"���9�I!��=� J�� �x�;�%B�h�
��K�r�L�X	Vl��.�pl�}5����{�d�SLޥ8�D�_L4���ݏx�=�YxF�@�%3͋�~�LJ� �� �����ug+]�@�Q8�R����-�ǻ��{X�Qj2K�#��qڙ�ց��}G��k0_p0C��:�xҍ1ҔE�o}[�+�O�&�pp��,�Cm<���ߦN���/;Y%�C�m�@���$�\Nٺ@*�a�6.)?	�����ۢ'6�2ҭ��U���Ǧ�>��X.ǐ@N���øq�J�ϩ�N<2ūɿ["^�5) �ś\�����G�������d����AVTp�^W(^�Q���.���1�����=/����������.�J���Xڵ(4'�\�Wsz�[%nV։��o��M�E��h}�ȤF��gX�F��d�<��(�/Lh2C	>%�����j�֬+�=W���
	x8��'y���כVF������%$4dZ�\�r�'����k�	�D�3�9;C�w���vzcP5�/��8l���Є��{֚K�~;��P�M���䎮+��k��LY�*�q �M��	MZ���jL�Q������ds3�8:f:%Q��"<OfNWH~���舓�·�#�m��Ϲ��p�VG�������n�{���ֽ����ԑ��W���9�p��8�R`;�^�ˆ�8j��A��Yk`�ꏪ�"���/�W�dO���ڢ���?7�}�Jd�GfyR��BG�{�c�%�� ?�l�U-�'6�$�5�P��P|y2_�����1xξ��;T����KW�����z��Nc��j�%j���/&
m7z<W��5 �� j��V��lyI���l��|�Ob/�5�K�0K�?U�G��C�(�pi2�9�� ���ixB$yq��n�a�#sxw�jd���h���b]B���p~Ǐ�ōOrgn��F�t�_�{��_X���ݚ��<����bI����RE$�2��,5�`C{��ʜ��X������|N������\>c�o�`�>�rf�u�� ���C�(�Gb�Dm�_�r�ALVt/���<�t4�����s��Ԣ��+��9=2o�����-%bF2~�DKsFRꠋ@l͎-7L���$.�xqGB��é3ֈ��'�V�v��ǖM
�o�]�\?V@���p.4���]EE�F9*�Y�)~0�5������0��tO������f��pg!��3� Ć�6��?��ۅ���}�������r��I���Bg�Nd�sa=��w�ԝV�[� ����A�W�N��L5�5�Ģ]��`p�%F`��ԂM��\�:`���Z��KG�F��rc���$c2��]UѨ �W�T�Ȧ�����R��� օD��Qdh'��K�b��5�(��7[��^(��o�M�$�D�g�%�s�N�kEj�W��"uAE$�]��/z���)N�i��F]*�1������>���Y (;m�Zq����`� 0IW�?h��O�"�_��!��@�@���B�i���\9
�v��Bʝ������]e%�	p#���~{�����@��W��������,��+��ݔFko��k�#w����S	�<ҧ�����ޢ��2�Dc[�\7Ku�gsTﶛ�G�JM�U�+�/{���H�J�Ed
2�$ס����g�on�GShH�JO�>b���}p!t8H�M]���oA�{7�;�=�/y^C��6�c�zծܗ>|�Cf�լ"0�j��������&�;HM��t~�����;�P�`�r"0G�5�4��ž/��sv����B#_�oy�6�!��^u8��X�J���YՔ�����w�z��������\*��.���T����K�o�����<� �='��/A�U��8k��惝�Pߡx�ᖥR�)&�؆�w��}w��$ދQ)�=��G��5	��;(�&�GI# V�OȞ��/)dNx��ǒ����s��قxM:�0�΍�o��5�jEp%�hO9�#[g��+�/ ��5�r��oG�y6�p�������,�j�{���\�-Q�����;;"62���S�I��^��P�~���إ�q�{��Z�5�=`����
]����m�
��1�ش� �9:�U)�w��R��WТ���� W���	��"X�E��Bpb?�X�͇����z��E����F?w��y���`�5��p��;��}R\+a$� �!F_n^E;z%�����5���B�U��N}p��O�lsߎu_"���?��( ��_1s��z�_�7�讲���U�ȕ�N��'4��#��6���N����$�'� �M/~���$o�5�1J���-��M�a��4wB��^wj�-�
җ����KE�ܻ��Lk.��.�i�߻�P�8;��M:��Ȏ��K�Q��TU[��OP�9�0�;�$4z��]N��A��6Q���/��;S��gD�mX4+S��f�q	�4#��j��[zƾ���}Y�Ga�so���Pү˸x�7�)�r��������`��r6����JgÁ�ӐEt�FC��Дj@���#�u˦3u�4M�ޥ�b���� ٔR���{��sXّ�Z�{K;���!%��Q�: w�}�$�����0����/�|����۵���6���4Wi�U�^Z�Lw��qb�?���g�J�	�0.�$3.A��5����EE��	 2�M�Y�B���F	����eZ{ss�ri���GĬH0Q��Չr�pc�|����R�H� �	��3sG��;��Z4����p�hD��sLPrڰZA28���@fI?S�%uK[S��oVȩ�9��VT-��e�!�M`<E��K��=fA�tv�K�v�?�����,�d7+@lxi���o��q�߭S��2�8������,�X���P�����<m��嘃����!X�U�_7G��b�����qҹ.����z����j��x\��M!-�.�����c@���1���H_&S0���˓���#^�R�R�Z��Ne�x�~r�J�#Lάw����^)]��d�н����߸�Y��=h!�;	�R���뫹Sb�!����g�1��Z�磞+��-�py�(1�)̼�w��\�F�
{|v������v�}�˭;�@�N@ơա�{�E`<�Ʌ8��#h�U%ї�e:M�|�i[���j����19�u1-Z�:+����&`/=�X�4V�e���-��c|`�6�|�A=�0Kv�D����.,���w&S�f��"`�	
14p���25����#LI0�?�D���!�^���y{F���l,��?Ӎk�p4�vqV��B�#��0u[�|��Ar[�����(ƌ������ҷ�(=/�rT�kŉ#V��z���PHm�H���j�r��yxkǒ~ð~!I��75a�+�n��U��U���Sj7�ɤM d>Yp����l-��=?_�0��R0���O%"v�@*O�b����IV-�ΰ������-E� /�T#0a�� ��D��G�5w�߸��wt�E��c4e�]!9����F���������F�bh �2ۻC���PV �bV:�Hwx_��T\��-}$(�U�k#	�YrYc��JrTz��;,��zpI�~��q�o��K���l��H��6#�/���~������'�E5tbW���).!���/i��!l��� ���8�آ�M����j�H=��B����뮄I\��8��i�f����E��>���]���ԫ����G��j�{৩���M�`�a�G(qO�`�{̬wU�cd�]J-8\�l/=-V�?�U*���VyK�<f�̩�ʩ各�_�H��w�-�m����u,�I�8cm8Fl���t� ^�' j��n��܏��c'Sx�;��I������ov�-����GQ��1_�g��l3��ͪ����&E�j�[�M��}y����Lv�ԕ[l so}#���ѯΰ�`Eg��q�����A�`6,\NǷ�{@��eκx'�P#1Oeo)S*�7�۳�$`v0AY)��W��������K��F�=	���Em'��z(]�q\y�wi�/ܖ{�s/Ҭ�v�g�,Ȧ��a]��V��Å�� D�K�'I��qa,G��������N�[����k�t��ε ��[��O~Ϝ�Wp��[*6�`p�_T�8$�HO���]/�5j�/�@o�LPaWN8g�PBQw�_U%�:��k�����П�UHU��j�T�뉵\:H8~w�2�;���+iE�����K�g����.�B�sm�NO}8��*�)��8ɹ��"��t�߽6c���ܣt{�t
�{&�����QY���eWOP�����v�ؙ$�V�ॎ'0��s٠�ˌP�:!�+|N��׽��3I�B����=5�y3�F�'F��>M���q|�����o�"b()�J�ž1������;p�Dg�X�d�>1��O��O�"�d)��/w��JBW�p���-���ϔ���Q���X�G!V y���r���;_�%�Ĭ
�8���G�u�uuu��
��ى��*�h ��*��+G���a�;�m���SfC�ux��5M�%5��e}�X��_������Rc�z�{�F%�ZQw�n�LmO��(�Te��En����:^����F-����~���ԹOV9���P���	.m�G=Dھq��G^y�!��r�sY`Q6\��(���{�fwݕL1���~B�3��_�Ծ�3C�Γ�a0���I(Nѷv�( ���~���*X��p���ǰx���P% DK�~x�bx��T�u%��B՛7��ʃ�Bݣ6݆,��n���&Zee���.��s�3e����'Fܛ�xՉ��l\�-.D�,���v�9�X��㲃�˺��#���1����]���.�n_'�}�7&�0��1�3�cđD�_ZF驃:>�3e�M�}C�o���O>���e����	?�&F�_Z�L��;b�7����r*����?��fG��ң&)_�%�ȐW��V¿{l��G���ʅ�դ7<V���uKaM���8�[����K�Wk%�oQʬ����C43st��JKy�՗�=�oQ����k��9N���>��Vʎ7�䎵A��Ezq�ЎOTK�F'�oJ��=l�~��(-�j��c�<��,�6ky��D���i�e�·)ء&�����L)y&�S$�Ԟk;�޵$U:��T�ɻ ڦ��j���U)sl)������9MC2X5��c�՘�:���j���d�dS�A���^L�|W[� �A&\NW�$� c(�M��1|��Ջ�.��*���A�qgJ�2��d�7�<�B@��2k�?/t-6MIU9���U4�OJ����2_yfC����W�â�˃?h�;�!���%��5>~�܌AAf��XΥ����fv������{W(wMڬ�4��xD��ɠ|�"��hĕ%�R;&����җ�e�����D�Q[uG	C0�p�}U.(%+���G���h�c�c.!������ƫ>¹^&S�ш�-��.�D�l`�tk�2���JYr�o�M7��>�*�Or���dE��4MR��E�:!�;�KӦ�ikq�������k�?�9� �.�^-���?
g������E�7k�dVex7�/�o#R�Cd�G��9����f�&|Ѷ�F��\k��u��7���֚��ƍ��sz�Ў������!��3�xf��4�|uǿ'}B���ҲwxBM�5��,C���6-o��	���A�&�#���?!�Q���w-(�/��H�K�	��$��Ҫs�`�K�:ţ+>j��f�^L�>&U��Yyo��Gi�(�DԒ�8 !��
�&wo(/b�"nLM��e��DQ[W��l�4-`I5[��K���ub�^�힛6)ycj�>��+�On��SQ�H&�w�y]�)c��U\��@H�	��@���@@?f?Vu�(<y%�F��_���$F[���<��	a�Z��',�F�2���d��#�A `�V9�9��BԀ�2Ơ����IX�Ϙ������
�H�(z%$�N�^�;\��Y�H_���j'@�sEg\s��@X�k�|M��׈��d����7����e �f9O �1bu*=��8"1����w���@�����7y���٣g�p�eo�ŰJ睸���B�9Hn1v����js4�m����������;#���)Ӏ��O�Ӫ@�A�XHC���� B�K�L��+l�J��.�����<.�ж�����4/ZIB�~!&c�e���X�I굙�w�M�A"����o�mtK�R�	���u�kC���q[j��neu�?3ù�J&���X�R�rC��pQ���e��tޯb1(Z��)���w-��z"(��+P�0k���ϵnd�gR��~�*<��u���
P,j;�_�@5�sa�#�4Sw1"�V� �v��4�?|��%��ֲ�NdJ@1�כ&��B������V��.1v(x�Q"�Z���<g�Q��U�6sCE	��NF(:���}�Jj�B�(��R0�k�X븠�G�-�o�FU:���e\y[	F_jA�.K�	���|�l�����R��k�$d��!����-(�Qu��/��g�9�&�b\���zu �s�r��o������&�33����մ�t��ug����l����������<�h#G#S���ڐr���˄�\W`2�7 N��#�ö��Ϙ������o��
K[vm�D�&t�k���Q��X��u\����E}����+��*�Tʂ�w߂�;!���fA�^w�K\�bjg�]�hɤ�V z!�M-��1�J��t���n�:��E�����
Y��H�h��;k@�B�"&Ry�� �ǖ�#�`M��,U�	�96�ej܏�������Vr�Ӝ�a.)�Y�62���NKS���j8��u��"~��ٻ�,F����cպ�Z/�}��$�ś�����\�j�U�����[���s@}|#�xZ~M�b�:P$�Ԗ�/��3��
���%b�^]:��E��W����hZ�e��M�9U��~z�����o�F�-:RΗ�����YkY���Z��.|����C�|���`�>�[ɲ�)�AF6,�ja��r�����w� +K���S��|����`gL���k.jfG�G�F 
�J�
����)�u-��zc?/=��U��u$i�;Ӗtᬳ�|&A���*�S�17$ZN���?c�2�����䂟sl/I፷���Z�Q�VRLdR?�}��>�$��d�����yl���ĝ�F�:�p�S��5]W��|0����,w��c�1����͞/�]|ӏH��ƻ������@�)C�ķ��׮�5LN��fp s9D�p���K	�����O����ӱ�9������I=�����AtK�_79���R��	�]X*��s+��zP��-����F� ���[B������ϗ���P�������"����.���}�����	�
A8r�<Y�C�4a���-ٳ+t���66U���&&ӣ�����4Y����/�s덑>�v쳌^�`���d�$�k��Ƒ�ቲY�N�E/KI��|i��h�Ô4�RFƠ�7�"�f�?F�P�� �7���\W�9�^����&�9_���ۊ�	�߄���u�V�IH��Vu�n�j�Ӗs�˽?��Þ��E�q�1le"���E7+=��'=0S�Ϻ���C��׈p+���%�+���/X7�%��*gc�O����T��j��c.�3�a	�PXq� �����R�܃��5�>9��&��=I'^�p�.�:*��BȞ	x �5^�O	�n1��p�w(tv{��l3���I���P�$�'��D*>�1,2!؊@�-/@&��C��K���	�0t�Ek|��?��Q����Q�2�jW�ӣS�.5�ڛH�������yt mQ)T�@�����Iz���x0��u�<݁��=q��n�ë9�|+�D>Ռ��@M��(e���(�b��(F)�R�8�r�܋�G�����7��~��N"���8��C��"�U
@4C�~r�8C5)^��4����.Ws3�Y�����9�V��iP/�ٻ�n�lt$�e�!��k��v,�$��4��ԣ,��Bow�0=AŬ���^��ºϭ�mQ�������!�;/�S)Ƿ�x���+i[�9~�3I3@²�U�z���?���F�s�z��ʑ���p��.Do�.;J%f8cO���D$/�;�^{g}f8�ZL�-�4�j�"��k�� �w?�~���ȳyfsSi���#��p;�� Hj���q�~���ّ�K���~?�> PJaA|˙6%t�1`����a�ڗF�#P����s�;;�C�ћ���TxB{\-k`��d-L�9(
	���K��j@HM^���i��8����YL��Z���5G+�"��BJ��"�EJ��&����W��h�g��E�!��l �5)+U��&+Ck=��(�R?�����f���e;�G���[5�v�W/�ӶgK~��0 +]z(GX�w��j,��c�3!���Dc #൮��%M�25��ոܡ�=�5�����;N?�����@����oi��k	]���҉J��X\"ǻ�0�����Vt�4U&��M8FlI8D�/�"ܦ�H`B�lU��]ll�!�_-]T�X�u>��
��q�;��b�^�v�<'����<���9�RXd�q���\�G�}���ڊR#:c/���^�\�G|��R���S��S��g? y�q�r���{()�� �#�7�x�(EQP�͔��W
u&��*8w���!2#>Q�km�#��kϕ,�>��2D��P�P^;[蚥m�6�?�%�"g�9�^Q�5��c��Z�|M������z��!(�L���;�璖��p�28�>�ט�	�B��!�I�)�Q|m:��+f�$�� o\F}&K΄z����5���)Յp�f��Yo����m�����ӵ�����*/w�]�F��2�+���2�0�@VJ���!�A�ۆ3��_�F��q'����1T6
|���N(3{$�ژS����I'?ݪ�6�XO���6~�{�?�+�} �c��P��;kpQ~G�O�F���X�3���p�q�rb�u�R/�����o��5����đ�É���-{u26��/�`�O��#FK�����F��k5+�=�����o�@o���V��9!2,S_�� �S�D;10�w>L�K�>�U#W�`p������N:�\�%ש��9�e2j���8?���,�JJ�M���9ū�l�O`�����7�zS������K������˧~ҁ�7�.�Go�]Y�������폽X��ƿ�Ǹ[TN���WY(�7�������L��^ MjA��InTY��FD��� ��?yC	��a�L�͠�����a7hs��NE}��1��#�s�J�zXt����=��9�����#���-��w��8�y�Q�5^��bDZ�)�,YS�yz$I�7��W�Y�y���M�rz�ޮ^���LM�,�Ao�fT^M���F�xy�;B ���8p?����[}w ��$܉34S�"�6#��&�^��Z� �ч���j��4x���] �f���h����y�0�F�CU"8��vrA\��J8�Z97�����	o)~��W?�����f�����e����z/�S���A�����''�V�$G�xX��Tp�Iy���Wh/�o=� ��� jz�.��V9٬�Hm�� /7����!N3O�jڏ���
L�wIt����377Y�T��M�ci���B��ｂ�D33O�vlY�g�[R����ύ���`��{Q찼��CcTZ�A�=Ѳ�ݽ��lY��0��j���rXzEߦ�ɋٟ0 ���i��UWܯ�R�+b�#_��]�ү���N^�r��P�{��a꽒[Z\@�Jћ�NJybgll~]u=bo$x�������z�Уke�����k��gs��0x��t�����UQ�;�ܣ��1�6.�P)�h#2��Z��|�!�@�ufQ�}�}2�2��)>����#(q����1�/K����8�Е��W�+o@.�ٶz���K)�&�!���$�7�ً,��F ��քˍz�PX�U�yG��h�P�N~	k;r�����Jm����[�4��d�4�K���VkW��d Ǖ�0c��8���mKS�� �y{�~���#bւ@�NJ{�ɵ���g��~f>u�#N�9��YW�P�l	�f����� ��/z�&.�z��8��lB�f�V�/f�v�3�,��G�xt4�3`��O�����#�SF����૊G���f^��s6&��%1c���X}�K�����k(�5�W�z$>=�J�4�������X8ئh��#ʭ�2*��Q��-�1r����Gp�!sG:޿���'6��p��1믛>��_�qSD�T�=!�`�cc��u?�ȹǟ�c��w�����>S���?*IC��2�F3��s�Nni�Y$�#���[J�����Ӹ�t����u7ݒ�sC7Q�m*:
��\So��R��tw.V4�N�8��9Q������*7�ǿ�ݷ#XVF]md@���m�/�;�:�~���[�{�0j�iѽ A�X3�&���ƽ��[h7G��r_�}�3�si��eWH�#���J9Uɼv��l8V(E�.UgU�L��U��n}����eע��	t���i)!�Q�t�XX���dH	j���Q(�)U r�����D�����<���0����r�S�()�*���@��U���ι�WQ$�.��PEE��	����[��h�J�K��g�KE��5��b*��r]�q+��a�"�[���|1Ij75�?� {���w���\��lù�	��W#��M��uT��\o�}�c!�A#�
����C,�6ga�\^_���t�z %��l����=�('��봃���a�56#gт���ﵦҍ-�D�R�WC�1�I���+�|��ǘ��o<v��ۨ�����1!Er��گIIwrNs� 5Y`�q��G蠀Ҽ3iA|��&m[考�c�L�����SH��UΌ���Nyo]me��_�t(����}M��8����3i]c�o�0W8_��U�w]&\}�I��` �B�d�����	�v�2F�C"�x�g�&p�)�~f[$�ƙ܌�s�%ڊ��.��_�����.���1��P��f)����Tb�%�2"<�
8.Un�0��\�ВXm����-v	߷���*�͐Mѽ��>Q���׆�u�I\��t �@�?k�"�㪍n���@Z����V�>�^k�0�>�%Rv�x����>�CUaIл���$9�lcz/�e�|�
�Q��ai���3�6�	ҧ���G� �g�!��}M�^�/����z��n�h�Hms��pL��T���<薏݃v�U�b�hL�T�m<A�Ҕ~Ft����6U�e��7���'g���L�y�yIw�d��P;ޒI�o����Eb��?W�*���0����`��ˤ���X��x��+Y�A1��WkLݗƯ��L��� @��-�>ڦ�rK�����6�oq?P����k���4�w �^�}#2j9G^�h�̔t���^�/�~m C��vT��;��&+}�q,\6V�V�I�H�c�Tr1O��-*���G�5��p'�
�6O}�:
iD� ��~5�%gL��?�TK^��sr���D6�W���t�������(6���5_�	X�={�#rǼ����7&���ج7{��� <�g�L!�'B�G�����t�k���?~u�7z(E�_#o�W7���������>��������t��玙3@!/W�f	�Hb�P �N�!��PBg�Ӣ5��k���(�h)��/R�X����N���p�/���P�s&�	���Et�Qz��< ��g�h.P�oh_R�5�[���p��+��fBAg��rz��qF�?�������xޠ����<�Ӱ��-��ǚ%�T�n�)�����&�,�����Hm��<�L�YW�U{<(<�Tߔn�(�����m`�Iqz�F�U�����q~~T�%Jw�"����V�Ώg1#��p���/<��!"��AY?!�R��_�3����e*��'�U�G':�XN ��SJt>%[��b��\�86�L1��Mjs вh�ZK��nҀ����`�h���2?wF���oψ�2=�W�m.���� �f����<?�� 35v\�����J��"L/�P�R;<�'���U�K���/����/���^
s��L�����r^��B_�5U�P���~V��7~6<.�B���a�|�8Yj��T��c��'��>�J��B��W.�`r@:,�Æ�.�a����������ܵ��9~v��Gm~���T��V�i`n�$���F��B�e�q��1-�- J]qK���G�K ]tԞKtSi�E�f@�h���$6m������٤�VQfR�֏���>�
�
0�f�q��^�q���a��G�Gu,��GD�2��s�o@Ϗ�A�2�!�:�_  H9���Q�|�o<��-:m�""OG�7| ��ޘy^B>ݚ�]�۹b�>s�~M*nE�l��ʵ��%�7s�k���R�L�8��~V"�4-��KÅ
�����E9������8�/N$�	����Bc��7�k�2b̦ �D�ʤ�]�&.�Yc�{}^9��Im���!,����oD.DT���T!as>u�gp� ���o�3����\?A4�Bsz�MR&�fJg���/��7���a��?Sv#�����lk�@�8BE��}��� Ms����:懊^�tO� ���cp��.\Q�����}�o7 ��ݸ�"�Y^�CҖ�l���Fy�n#Ȉy� �`���Z�8u�ca-�cUz�������z`��y�y�����Ff���� __�p�qR�f4�ԉ�G3�-D���O��',� �4�?>`}���!E_@� �s�5t2*3�w"��V!�� �'F��')8������3� QMT�;7~~^�����YγCA^�����s� ��]�#vm�K^oS(��<�]��"��0�y̖1 ��xz���q��{4�գ�T�tsX����{� �&M�8���3N�~��Hr�ql�CC���<�S���h)T0��W�WVD3
�Y�>E��H����ˣɌ�b�£�������;!�7��0]�rs����(�`����>�Q�(]�!�w��̅�d�j콼8�Y����jIЌvtސs8X�8�un�N� !w���[XҴ��oF��߇��+ur�C�<q1�q��ۆ����0g��Q
�˞��4n��UpJ,�<�f=���"�S6�w�5�"s�O�"{���Q��Z�u��'~�(eD���d'bְl�:[l��4OhP���N�~�=Ǿ��L�_,��5Ūo�f�g$ut �
�f�����'�ʂ���M���,�Φ�2�b�Y��,Ip���em2o@�j�� q��>�I9�*���|��:��O��d��ߑ͔��D��<���J�D|��P�@v��.�j0��$��s< Q��(3�;�^�v昷�Zb�w ?�Pc�}#��Ƥ��As���:l)�\�u���Є����|����~V��o�20J��7��B:�d��ʹX9�?.�<e��~��m\	�p�k��.��$� Vk�5T �SF�n�l�lǰ�	N�v�: M|}�D��](�N8�=ݖ�W)��d�1}23B����2�c�9��̶����B���l��B�� �S�h[���~����v�CzZ���B$��E����FGJyl�)w��#���{p��t�E/���=�)Jl�g���^�i�4�-��N�4-ݴ%n��C��`����"ڸ&R?�tt��U#��⫘�'|�i����{��@X�ƺ�=j�@���0��u5�����%�7b�Kw�ߝ�Ϛ6�ĮA���L�&1�=�%txY0�vN���5{k.+-�:Z�8���20��ل&ÌU�4�y��ۤP^C�"���ݠǙ���
#��T����xbn�pt�X�R��x�����)��k&�\�G/��[t�?(�8�Fg?�(�4;?���r9�o�eǬ�*pF����I��(`/?��0��r�`��cרo�z� �����k��P�i�i1�v�l{�[�9Fx�$��N��3Fy�U��𬟶݂-�����VI�l%���6C �
Yj���}ܔf�q�X��rN��ȫq%��_�se����i{Hv���IwE.�k3����!<���)|�I��V~�!a�U�W�ye�Hr9���{�uLd�ɰ!J)͌\ �~� *{�YF����X�τ{M�e(�2�5M��~]-oJQY�L��C)��ʜ�[�d&����X�=��
�[$e�\lZ��
�F�˗ZXp.�yU����$�|	b!���Bp��nb��1�m�٧藵����5�0�/�'��U���&Q��`�(�T,݇l��|f +Ed�0���lV��eB�z�|�9�:��ʋ	�VW?`�nҏt���Kfp:�G�@v���:�h79�l�Dg��6u\�<����J��;��g<��t��
�T�JΫ��Ez+���������7�X�Ǜu�25��$i�	g0X�=�5X-���χPea�J,߲��'�~<�3EC��tm �dZ�ZL) ~D����P���#�ĵ������D�^�$i��-t�+�4�,!�T�%���"�f�>G@�7��ol�=: '^q�� Mk�wY�A1���7�%|xM�Q���k��E
Y�1nǮ�	��}���$A����@-�O��:O_6թ�̀��������bn$¼E�<.f;��D/$��跾�W��`�e����^ �F���z��c���fJi��_�=���>nEwG�"����S���V���?��,��vXFlM�9�^��gb	���X�*���6Na���hV�',��(SQ
9�.by�Լ�N�+J��X��~��&Y����_b�};FTs	v�t"i�#g�}4��v�x�Gt��T�U��_y;nUF�7*^�@���@\��x�R����\�0�l�,
�ZE�J׋�&VNP��wk�� .�_�m+
��"�F�Z%��2��}k�$_�%�f�r�Zi� �;G����nO�D'�DQ���B7r�!������6M_�n#�7�$V��<�F�Et��pr^�w"*���h�������_��]V��$�^��e�y��S��@�	ŏ��I�^�����J�0��BO~[Nr��(tH|W b!�J�����6��C�=��(�L�K�;���g�9��o��$d��8��vc��$�QWm���@�f�鮳�İ`p�=�@��QaИ�l�]���8���6=O$mq�X%�/��	�.?Ҕ�HK��	�5�O��� �JD���h��zl�~%+i8��.�����\�f�.��0��嵃"�y��4<��I��ňζn��djl�d����ꂬ�&�,�����jp���QQT*� w�6JYֆ��j(�]���Ki���V�<�����No��wU�rt�����]Շ�}x}~0�i�ǉA(Wi�Ő�����"����-ÛvH���a��{@.��W������^���K�%JS��{���;/Qh%z�x�Y�x�}D�{/]�Z4��C�L4_%���0�`U�aSj7v�vI���nG�H�3��{��[[�������� R1�j0�ft���&�Qnn�Z�iV���]��̢�сV�H�V�G�K*& �y��z0*��;�H9�^6���U��W�����b���YO׶�w3;�W�Ê��'TJ���ID-�)˺���z����J7���Ѓ��x-��7�V���{�{���)�˷O]�<�0�y_�n�D}���UU����,�iy~c�R�Z�Nm2�yz� 2�:%����q��hB��i M�����un��p�))Ds	c���EC�VM�N=�N�
��#Μ�	_-�懴�|sp��2{Uux�MC��*c��p��������@��A<�bjc�cEd,�a�N�IQ����L�ǲa&��[�t���4z,��P���,q	������U�^��:>�5}���MV��+�*P��϶T޺��r	�xb��:�)WZ9]I0P�!�[����Qk�d�C!���k#����k���nՠYI=�b7��ê1k��^�
F�����u��j�x5݀J��w0����J,�B��d%��c��(r�iQ�VG�:��bI��A@VY�����7М������ \FFѦ���ȣ̖�gʭz#�o �$���F��tY@����Eş�-[��m\�����okt�Ls�]k�슑��wgD��Z�[�Y�_k�m9l�J
�M���>��SJ��<<�8v�3ꅞn����Y���F��s�w���P]�_(���g�S��-�g��>4��.��+SG��j0�1�C��C�))ʒ��R|R+Y����;P�׾V�$�D{�<�nꃿ!) sL�Z�D����$T3�1��� ���/�mw
�������cҼ�G�a�!߾0�~%{̹�p�����0��������Pd����CF���E�Χ��0oi�(;�;`�N���
�?W�����E��D�mw�[��E,Zk|��VL��>�Y*5_�Ʉ�,w(�Y������@�7[5�'�����xՑ��c-p�f!�;F ����D�E�C9{9��?OGAD4��OE@``]u�s�|���q���ObG剑�z�P#��mC8��ӊ��<�G�)�YXf�g�o�7���/�ª/r�jyI�?�l� ؼ����s}q1'o��0���j��v���
��5���o-���E$���cЈ��O;�\3�6㢞ZL�F;A|��P��v[���y�
�S�8�}�i��L';Sn�}(�G}GG3�a�u0��/����(�t^E
X�65�Y@�3�-s��ukML)\�� �z(�9;��k�:�H\P@����˧rQ��nT�=����q�� b Ew��f�&U��'�D�t����ԗd��eTTL�25/;�ƵD�Y"`�_�x��?��_������Wk,�C�U,�@*������R��<�_�L��}[��V��_V������ai7�\���s-G��d,��Y=�|�*rjsG�oPoB���=�C�1]�7o��G�ݫwalȺ�Ey'6s����r �i��f�_h�Yw�m����۹"b)��u�������i"'����Kj�~�����+d9����9�x��	�M����l@�g5b�O�
be���U��A��@#J��\R�x�ՀV�F��8݀�－��Ra����P$R���ب���>��nӂ�a��'�� (�����^`_$zж��}�G�Pjt_);Ж) �O���+nID�1w�����(���˿��ؕT+����^�	�˓퓙=U��)�L�%G�������hW=����/M�%~v�n��Y�W�C5^�Xt}�)>Z�x�� u��\` ��+���֝���o�uU� ��ޛ;@j��74�[�?D�]�,��=��i�xT��z�t�'6���L�?e2� �yfz&�I���?N��\����t�Qm�M5���.O(W��zћ�^�\mWq���Fۀ[�rGlpʇَP�/���M�z�-�i�J��ԗj&����C��T�1'�t7xJ*��;�?N6��0�q��V���c�0�w��Vjӟ#dg�`��75MK+V����ى�"^�1K,���!ĵ�V�mh���\��+,�;u Ѽ�1�G�tI^ͧ�>E��m���)���İj��3���g�a�.�G��n�}��岝�|WQ��{��oy��/3!#U��G�y�/�I6q��!���m����gVyUT�r��8GQ��5�O �x��!�"�A�$����3��e" U��w�>�	���B\ฦj��2K��.uup��H/+���X��Q/�hNsD@��� h����S������=��X{EA$�Pu�5 O8�!|8t0ѧ+���K�J�����;q�W� �Ñ���� �gϖ�I=Qe~2�[�N}�c\���-n.̶�5�-�{	/l��� ���b��?����B���5N� Q�G�m�ӣ0؃#1���<a(&MWlS��ts�`��K�[�E�Xd� ���"��DKU]^ =��'�
f2;���&b���C�7�+#q���(E�� u���O� Rl�7��4����w�f����¦����i��UA����c�	~��'nz�| m�y4��F��FJ*�����F�}s��9�n����$>c�}����!��d�ҨPM�h���c]ny7��kޘ<���3�C[��P����k[�����쥥�8�B��0i�G/�`�����S戣�~�y߷py���q�����Ɯ�Bo1�-h$� ��-!�l_R���Cg�د�2�<IG�X]�ɀ�Q�ri���8th?��@��R���.���-Ohc�?���_�3�y�|̞R�_M��+����e�ŋ;Ͼ��-Z��g�#������_؃ˏ"+W����h(L���������N����L�H�3�p�uͷ�SvxBQa����ӟ�����Ez��_��U�W�?N>�M��r����Ĭ9�E��%��������D��Gu<,����n�QCa�n�݂�\�"G�&P�9��M
�3�Su���fe�� ��lTS7b�g�?�|]<?k�T�^�Ջ������:�H��ϔ�4VZ	���
*�'�2j�f�g	�#�>	����s��$>Ҿ&�����߿�����^C���2P-P�C�ɠ0'�o�K
q�y�]�/��G{��Z^�_�~������>��4�JCa�7�^��i5���=�������MR`D�?ӀPH��g��K�ޠ��Nc��c��N��;�}�u󎴕���K��e�r����3ܭ��_7��u3K�	πRw
�]�B�ݾ�(�������X��0+�7�0�����B�=��3V��Ԑ���H�>�E�������r���U-���i������M�< \�p�!�������~���[�&��VY���A�}(Ӽq٢�����y������_{����[��u�;���}��`��NA=����ٿ�������G}��_G)y��U��{|BQ�k�K����"Jj�4���#Gr�3�%*���ڔ�(֠pǱ�x�\C�0���n#͓\��X�hl��|��f`����Ň�
X��G#��ݢL���m�T�� �S�⧰ǡ�mϢ�5<�a�M�E��ptP��;?�M-+V3K*#eO��s��:��_]�nA�q�Kv
$� �G|2��|�Or	�'>�6 ��2�˼r�ca	r��4>ܶ���l�v�Φ=<��HW���
���q����}
�8+��6(B������L�r$t��KN_��Fq9�����]���6Mo��)d�&{
(���8�{o7){(3��e,�`f�=�RI�J<(-�ק��I����NM�Wq6�5�����i)��zw��}� ��) ���V��qr�RM3�A��pm��Q�Q��N���(�K��|Xpcg��)��p��}��kgλj�X�BC���[���a�M�rSjl)�Z��g��������bQ<p�G 1,�t%��~c@�7�S��[>IY �����VΙ��(���h?u���J����� �u�%�)�8X?��uTG��vL��@�&��G/+�i���q���sR���,�[�h�<Z=�y��|����,�$OC���m%�t5ì�XՕge��VygI��rJ��
8�N�AW��L@����{H�P�����qXv�,�ΪB��,��X��moDlb3a�#�	�js}�J��=�!��IS�q�Z��jq�G�c j�Q�ҳ�"�ݮ���k͡��Y3�+X�3o]b�2w������"�� g��dz^���+�7�l��z���ʚ������Q�� �C�ID��&I��m#"�u6�����Ȣ� �T��[5��^=��7�M�<�����l����1�7�M&Y>M��[m��#*�����武q�a��XC���(��A��H��N�ԙ�5+Љ���b�����#'d�q=(�=���Aǎr��gL��}��ƺ�� �|��~e��X��v
��z�\�c��$[-Xf���y���}n��	�ӭ������~C!�5	�7_�
�������-C_�����$�<��
_KYs�@Wm�+NYbI&�a8L�Q@�m<`��,�GK�J$������
˰/_8-Kt�ʑ!�Y"�-��5!���S!c��f(/��j'Q.���r����#{��ޱ�xԳ|�����R�.���ڻp�=N-}d�^�B䰄�	� �5᷏O��8�4����B0cE���`��3��hoE�;e����x��ݓ�F�����/��0��S�]���!�34i��u�<��,G�s�m�G(���y)V�K��߷���Jv�
�
��xW(�!����_��@��6B=bE���.����(i~�R�kh-a��1�{ּ���&��!ٛ=��k~fg�D~uGH�fY%� t�x�C�ݫT�Tʺ�ܶ��GP�Ki�N�
Gjw�����ag�a�b�'RX��y��&�_��W�>8p2HV���Q�"s���-ǅo��C�#��W'�qQPv��~;���6�pW-�c�T7��VV3E��]��v|vy�Ek�����u�$'$K��ܑ���*����hө��&#������j�oimH[	�l�+B��˧2��I�%z['H� �.5y����hR���*(M=��wol��m��J��K���Ô�DBa}�3D�H����!�4�e��_dFK	�3�J�>�D�D���Ca����b�5V:�Ml`a������⡽Ӭ��03?9DRMr>�X\s*��:6)�����A\�n� �(ZC��㋍N�
ט�ŧ��<��Т�&Ӄ���E2'���>��s8��oF��x5����.ݔ+t�k�"�X��ӅZ�Fq<t�����aS�V��ɴ7�UT��ke�S�G߸F��s<>�]S�Ȅ��_0�� �>)�{��ny�L�j�	(�)�ؕ�V��{�P��x:�>1ګk/@Z����ۛ�ʘ�!�8y�''���	���G�~�M,�Ч�eh�Wқ1(�Y�&8K�MM� ���\���Ḋb��J�������'��:׋v@�aD�AN	���t?x^Ke0z�~I���l��	v�|곻I�>�U�D�v���!6z��U����P��ly$�F;P���7�zI��+H�P���p��ta�Ds�G���v�6�.���G�?��ü�Z.*l;͗~?9]�cE�t��)�&����b���u�>�E*"R�#Yc�Ma=Y�V�~	��8��>�����SQwƭ��&?K���ޮޞ���<'��t���9D��n�tlՉ�[��SM�o۽r�,Ө3r�����*ws������4�����:3g�{�QF�C�M��ٿQQ���7�7Q@`�?�	�Byd���e��/w��i�]@/�rm�]΢�[�%C���sU�V���0]���'$X���g;�~,����D��L�݈�/��h
��-� =+3���}X�Eƫ2T���3��3"&yo�7[����7��2��瀀SҲ��U�eIg@�Vfej�c��UOa\�t��h�Fe:��]-O����ٽd�	tVC-e���18g���FkUCn������ϖ��j�z����u(X�"1/{�����E~��3�83R�čZv��%�(>`�q#�+��-%܆�>�1���ſ.�G��3����;s$�EO�*A�J���#r3�v�4s�r��%X�z,?��)�}���ÿG�A�0��2�:�9We����E~��R���+8Alp����Ϲ������t����~��گ�&Ĉl�n��:�Z�U���a��/���)�h��b#P�����"��8.L��z���z�~������b-�F����8b��������T�yܴ>6���O���z(�l"�	|K"�.�d�֏���@ƂF�����1?���-F�*�h��;� �8��ˋT�)���v�sd����LL5�Z�Nf�zz�aV�
���O�
uA)�漇K���{AZ�y���|%*�N4�pg����0�0Ψ`��q��B+�w��Ug�O�7-Jq��J�u��'��~?3���-תR�<S�(7¥a�	Ŧ��m�m��+}SeQ�6?c6F���Kv03�n<s�Zܙ��[f�i5��4��_m�n�˲-�3��Ѵ�D��ER'�:p�����A�lo���-�&�o����87����
��f��U�(��V�*;��0(&!a�l"|�+ޠ�-9a�D�$�+�G#�[�R����uM�IW�ii����<�c)��*W�Q�E�W��r��>{�����p�0��K���°��r�@�[j����,���G�T+������Ns	&ۚ?o��U��`x��l�F���	Og���������6��}�2<��v`q5,�'WT�j1a�ۥ5D;���"��'���/��	&$�#n����eu��Ԙ,A�8o�ΘCO41���^1]j��J��{�5)���������}��A� ��2U���It���۳�J��ڢ�xrո�w�u{�(}L7�����`��h���i]xݱ�x��Sb�Т�V�c�,�9;8�V�X6� �nҳh�qt�Bx�2����99W�����!�Q�|�!�(�ܸ��t�7 ����dz� ��{DT�I?�S9���, �j|���j��;��m1�1x��2xōs1q�.kh}�ׂ�_������ɯ��󑉊%���}��W�Pה�l��@IbI���j\����S�@��ZV t� }r�6zέVw���%��*���Pɲuh-��;cI��jZ�)�N���::'N&R��˷_����}�FQ�,���bB��?�� �1	�! q���BqY���=F<ػt���g�L�؏�{�ފO0C~�^�	�`4	w����O�_�.�bo�yW�}ө4&�g��j9GG����fL���3R��YMs�#S������ !���W��4?��w3��@,4-�Eu�] �?�3�!Ԣ��Nr���x�f���;�޷D�{k<�e���w�e @T���K���ehR�`gO�ո�o��˾�E�A##:�X1Y��z�o�Hj\�/T�_��r����u�0ֹ�n�J"���0�ӹ��WA;�Oiy�J�G�#l�y�/ঋ4�;.cd���v��,y�};��j�k�����b�}��vt��~�y�=�p	�ﳛ���p�N����3Y�������*���k�O����#{B��*c��6�s�a�A^m��y�H�ߔ����Q����`�,؝�y���IPp4s=�V��L�D��:='�C�ei� �)?ߎ��+�b�������$�Ц{)?�h�o�M~ogl's��}����k���rZo��|!���t/�(E#�D�I<����(�"��v�b
���Fa^�I'�&�g�Ї($@	����w�I],��Q��c���n��ɪP� a�XutLdD��V�J!�LqHdc+�H��T�����sG�K�3Ϊh%��٥gIJ��3u3a�y����{�g{��
�I=��|Wu�&���bte9�n��,_��bJ��eXb��!�$��rF�f�b[9���1�s�� �8�ST��������v�g5����_b�mpj�8a�"ֽs�{�-A�\��WE �6�T��=גrĮ)�j�[4���M���c<R����V�B����nF<��� #X�D�p�:J5�����6����~�F�_������Eppsݓ&Š�����]�%�f���i|,<��I���"�P`�L���2���Z0QX�X9���~���:����H륓%���@�t���9|֜?y$�����V9��[p�2�iW_D���08�9��m5��|�J�c&ef�=w	�����Z�BL��Ŧ��(�V�Z��z�s��]��Rcj��fh�T+�x��tY�IM(�fl�k����1`m����-�wƧV��D}�c�HJ���)>e �9�����S���9�ҁ��2�"�hN���~X��;E�ߋ#�
'0u�<�4m>�f���9)�[��쌡���H�[{��o@���P��:�W�k.�*@�WS��P�7�,sd�?Ա��5*���ƻ{�`��ӻ/�~��=����qv2Ӟ�i]D��[����By��m��� ��ߛ*揋t堫.s�&�kJ{�3���"�����9�ܬ����-���~�b����Џ�U����\�J[RQ��	+Z�Y��M��}ٔWS�{B�L���5��ٓ��uc�v��4͚�86p���S}VQ߹	iK�B�N�3�1�_��/��������+�k������!Q*$�R+Г��#���t	���}|�d�Q%5��X \��͞]qO��IJ�9�i��Ϲ���|N�6{�F lSK�;*�����qm6&�=�K�tU��!��!,RW*���9G(�޷�%�o��!J�)���հJE�,�! �������Fx�DK����B3�����A�����灿���J��a��Ŝ��z���w��,ܽQ���뇛��t��U>�h����)M��ܖ^D�5�;}=x0��d�ܫȐ��qT�$�5Q9��B��&<E>�F�����g��~���=�Nfc}������pb��	lD���2�9�g:h���-�L��^t^�B�V�O<�ݠ �S�eX?xO�u&���I�UNG�ۭ��r�Y��xWS�-��(µ��@	T�z1�.v����(�B��x��8+)g����e�p�I������&�԰� BI�8� r�b�{^S ��@?�����\�q�"P����g�i�=���U�(�)�V����p�Ks�����K��$�0�ח�j��X��.��@h�S|"Zη��z�tx{Ďa��i�e=7�z�wpƏZ {��s���}�+򇶈R�?Y2f�Q�O#o���LJAK�Z��Jpb[�.9���]k/�
���P�L�)���m ��kj1��'M��D�?1����*�^ <C�uW2�TDX���",��s���{Чrp�FZ�L��y�k�uL*�&ǁCd'�"�^�2iL��q�?n�)T�ے��&���/�۔���F�<r�RN"|saM4��5kɆ��FEׁ�v��tu�J�[h��B��H&+�<�����KQ��s��
A��]�y����<�/n���?8X+��T蕶�i�EI��.����g�Z�Ye�U͑Ɛh�^]�,4����Ck��O��ВԲ��37W��^�6J�^�q��+x��.;3���\�~(Xd<�+�"�O��S���f
8���T��O<|t$M����|fn��8�g9�2
��}��02��&���U��䮁P�e�,J�ǔF�h�ݍ�u��������9����\/F/�ZFHZ	1x�^���n��̥�On�#�3\hq1��$5� ���S�.ksЧ�r���b���j��lLx5n?-و7 I�qA�-�tZ ��[ɾ;-%!G�n�?q��d�I?#Nj�m�F�q�UR��	�s툂�DI���{]��&/W��W�:�G5��|�����]7[fDII�̧�j����R��2�"21,����F�k���KZ���bl�6�k�� u�o'bxܜv�N(�+Q c'C��P�������{x`Hj˔�,�kŏ��5<8}��oak�<���i(��M�"��� �'�o6�O^�� �Nr-�zj��±�5��!�+/PR�6�I;��Қz���K�����>A��Nwmd+k@�[}�Ƃg��ܙ��V�ܺ�N�4��%ԞC���*�-1T΢�>���h:R�ܩ�N��<�e�:O��S���� ,�W����:����IG�0�Gs�?��ϯ���+a✍N&���\.�2嚉_%���~�%8r^i��}�` 	X����Ↄ��[H����r5]�o��y�ɶӚd/�	��� nV\"�CE{0eb��� =;������u%ݡߚ� ��Z-'�2�?c��%x6'�!imn����exP�����e�(�f�c�0͟9Q��~V,�c
��tB��ډ͍ޯ`s�Tz>
��Z��,�� ��ym���Q���~�yMS�1���Z�w�
tR�Qh���]cl����Dm�P��1TeX��K՟��R<f��!sLDt�� je���~�P�{�j��E���C=EZb�n���-=T�k}���@fK����[�F*.�֞�F��)/n�"<�oa�K��<� P@a�c<��@-f�3�ЇƸ�8��$&ʀ��0�Gq��"�Ee6��[2�<J]�"Nj�E�P�g�!8F�����l\4�аG�����^`d�_�6d��¯�PDX9�d�3�Ӊ���T�ߌ�D��o�@�q����a ��:Ͻa����:��`����	F����ֹ�9���}�_j^\�97|�pJ[~���,Jx�E/E�<�0�:*X6�aޫ<}~�b	�j3��2�/JG�ئ�j$���{S��cu9�uN�S�f��hC<T9��C,��$��VS�w���33��t�la�
?j�%�VJ�Մ�^&�s��0��A�����Ӑ�^�(����y��E��Y���cix)v(6��fi~��#��S��E����Ǣ"�=���`ނ�p��lt��[^�w'�C�vm,�=�����5*�Ҥ���C�e����E��n�B�A[!�����=b
P.B����3�T�>�:�X���j���{{B��@Q�B�At���{t"�����nv�`�����1��/��~eH[QH^����]�����,���c`�4��A���-d��Yw��=�2�װ?�Z�'�{���c�Ю��n ��B�{�iő�?�D�=����J�54j�4،����!`�j/��Zc̰	g+��?-�eўJD����c��	Q#r�H�g�V�%À���,S��J�[���l&�B�sw����T�`t��B�v@"^��s�\=#����.���o�f��(��_L�)/	�׶�PM��������.���+=RmOP_Q��2��*�_����qF�'xs�F�x0w� a�Y��/�z��p��pL1�ugH����e�l�O,K��h���{��*�=U��G���]��a���8��z�'�5�Lpo��P��3���>qm(X�n�
8&��P���H��Q���*���4+� !�#�RR��-��i��}�1m�79�%-�Mu	�6�j{�0'% ��M�Z��>8��N2�m+㵫<��ʥ�M���Q����.���ۈH�
W&���~�="6K<X�8m�Y) S�ٌ��Ə4�;��A_=�C���� U+]���(}j��ha$��ܫ��~y	�����$@j�o'�hQ`��.��# ���F�$@G/���fR�Ҥ]&����f��#x���Ge����B`��
g�FBh���ҰV�[�D��R�;�MBy�1X\{��Q�3�*�3�V)3_}!޻ҵ�i��U�^+�>�����f+���������%i�j��L+.��4$�@�9F�g刍K��C�3NM�5k�gՔĺ-"ɾ94����s�in%�;5�VZ�=���}�����2�d9w��_�'��X���YO��Bم�eCwYD��v��'��OTj.��ƏDT )��y�m���=�>�Go-!}Q���2jح�S��ՏA� p���N.���⥦�d��?t�4�ʃQ8�/�@O����)�v}�M8)��U:�[��R�Ζ�+N��9�-\0�3��G����Vu� Oq�n"�$�#b��9ͷR/*a�b����H"��������ޔ�OH�HB���z�rK��mTU�	��߬W�@_���D܅��%���)��2hI�L[�ñE�{SE:��6f�[��J�t��l\d;!�YQ�GhK� �sդOs!��\� KsYfn�3_�C��9E�G)"�Ӡg϶Ӭ�QwA.j��l��D�O����Ƹ�)��.;#�Ёia���Qd����=s\�~��]���}�W���F�+�� Fw���q�����v]�WiGI��9��_{B��3@1�^~��w ��)lc���zDHV#P/|��&�\��2�=s�����e__dj�XR1�:}_&����j9���çZ�ՌT~����9fS�>�ty�H�ڸ�G;vfƟs�<���#|�5Y�O�B��v	�Fs�I@�wP�ln�N%;���A�l�zt$��RHZ�z-����]�Ps>�4���i�yRK��i��D!H���}P��ى���J��$w�,��M�?8�M?�|��߬εL��Ln��uJ[�#�oB�N���)��BSX6��w���l�V��p�`1c�:^�M|�gs �������̟Kk�*YI�\T ��qW��!�c�?�	�x�`��+�R�&�a��*�K��(Lv���C�K��ؠ��z%�f"�_�O�� @���Wپ���zo����$��&/������o�E�	�*~-�[0���2�C���^�qu]���Ug��,"���=:>G�2a	P����E`�'��!$�섬��c�R�W���ĳ�`_���r��k�P��d��CQ�]�%K�k���oaC��~EٔSx71�Z�����JcLȸ,��2�v���,~V��P���{W�x"����Z�Kq;?�_���v��&^��tԷ4��]Qk9�z��NZ�=���>�p��8$ּ������@n�5�p��}4����]�Z�L%���47# �̄��_�j#��� �[�je�n�<��s�U���C⧀���	��ǧ~k��t��{<t�D'��N�	OJ��o�)����ٽ�;I?�����5���,ϵ��]MN����>K�O��O�n���."��(�Q��-�NnE$�4��Xً�?ʜ�`�?	�D+�@@��~�3Ԍ��*��]�6��!�Xɰ[�z�	��Fk�N6�����Y�9-8Qn[��6�yA���S��]Z����<�>��Y�p����]컂*|�&?� �MqNd��1iH'�&�P�^ǋRv\b��g�e���7�(y�d�2�����}_�PP�V�V�PP!��OX�_",p:3��}s>�dv�6΀���=P�Pox{�2ƶ�,�����|�fX�us�4Z���l� Zvp�JM�R)�Em�f�#-ݼB��Esn��1�g� ͆�M��� ��{��a6|�x��>�HT�$��q�Nq~�� ]�5�֧�PAG+nؗf����O�v{�{��@���.�K���O��GP	�OUr�& m���8��ǵQ���sޜ���S.�c��x`]^d���*��?��㖨+�c�o����Gsp��ҁ�4�+�7��O��!�<.�l�KP+�@aos0�7#��d'+�&J
��mX�Oqi+�Ax6zs=0�������#$0����?�3��ɘQ����.�H	t�
T��3v�W�i�j�bzD�G��~7�V������#�%��	�\]�~�%�����eԒ����T���PY�`G�#�HO�{sz�G��n�q��Ʀ�SF%c,��q����!�W����@�6���;�Jh�^��SK�U�+M���	����FUi 
G�������D�3P92�S���Z/5a�HaP����E���#�~
c� �,g�U;b/�?�qD�&�au!��;��ʩ?)�F�UO�Z�0�)u��0�*���k��mI�X�.T�>���n�뀠C�n�)�
^XCKa�tՠ��?��6a����8�i��L�c��t�^�t�-�L5��Y�T�AoZ��r.櫊���S�A�iV���k2�D ��r/�1�o��1���^��۲&v��Q��[����U�D�Y�/�"eLkq�
�d_��\!*Oȇ	We_�yH	���/ҍ)���$xO{E�x�5�5�s��(�3�F��k?�h:�f���:��$�q�\���C�o��y��ɋ�O;�㗹�T��,���<ї0t�C��M��7ܒ����s#��Y{n����uJv�V�b鼉�[�~���x���x.�>Y�X�Q�*��=B�u�$P��DzE����e�(A�¤[l5Ȟ�:V�yv�,a�̓T.)���o��T,�-4�8��vb�`������'HAW�SH#Im x����� :e���/���h��*��M�Cd��i�*�½p˨�i�)r���R���d��`���'�{P��2s���ȱ��E�/�����������
`ݝ����M�`��P��X��r]�GТ��M���]A��u��Ӂ���!K�2:�!��I�b6���TF�ObӪ�p�'�)T�c�D�8��@��G}�O� ���4l£ysr��'}��j�Rfxۥ>�ّ�;d���C�y�4,dl ���*XroѴ�4�4'K(F���:�A�� ���S\&!�{m+W�?l�ꦑ(��02	�Q�b+�&wh	�^�\t���`a����^����ְ�z�&�b],yt+�Le_3�������No��%�yn� ȷ0�R�M���wM�1��7�f.��wI������m����+�o�|ٙ�&V��	M��6�V!n�>ᓰ�ǭ�ڙO>+��T� ,`���1������B%+oH�o�8���.�6���u��$�y4Ȉ���=��7��ŇX�0��ɲ�'͜G��;�CeqpZkL4]�_�B�'.94����\�I���mc�_��-��~��.1~^+KR��i����xBlC�h8X���g�Q����K��mv�-������<��N�pK�h|тHF��GYZ��cJ]��l˸�D�4vr�=6]x�.�Щ`qL���_]��w��� ���~����fxes�G\�/�_�u�̻��%0�wd�U��J��;��/+$�f^��t�:�{p��@�C����b�$N��ɗ�Ӡ]�b畚2'����sc��0B_r����PB�}�:. ���c�q	��Y�񰷠2d���N��8�)>sj�I��#K��UD�.�4�`��3j��D�v�N�~B>�J,������ CVB���>�v5�_�`s�F�\T��@S��#o���������%�BZV��G]V-��5�8u�R����1�u��8^/�v���ՋQ	k'��_C�| Ւ�\S�{��N ��.\��k���N-!��#��l���dGȞ�}�Ow�e�4�_L1��멶B��I��G2��B˷�9J�[2b�s���z]���'Xe�L���U?ܧ���|K"�1��q;�����X�&�~o�q܀�8��A$�j<��S�b/�T�{+w�B +����e9;\����`pÙ=vŢct�j 6]��W
�K��t��h:�:�:�g���_]��\ֹov�$�#Vw	x��-�܉|)�*�0��9�"n��u"�C_��nU���#�W#� ��ؙP���vU%Z�(�^Ɂ\�ȗ�-R?�S"V�r7LN�P,6N��ЀI�x��=�����hc[z�����<��S	舘�YC�K�3�o��а�����
vo�W�]�����j��k��2�L�t������+�젗K-U.���AP�8c*�Ⴈ.v�d�&/9�1�u���!#?og�PMR�?S��Nø��њ�NJ_>�(��oc	dw!'ф�r�L�u�FS(�>nl�3?>{	�A{���ܘՐZ����Zw��	T���}ҭ�w/0L�e����)S3���7DU'�>o��Q9�[����BK�2�L�V�YʅxM�[|����u����.�PU+{o�������[���G%bL[�Q�h��-��\�j6R�נNgFMI�$�<��)�o"`g�IԐ�Sp��l�]a���f��ưq�(e:��ŉ�̩tu��j}&��	���<j���f5�ډ�@�� Hm��c���i�ɸ������Y�P�/�����
��]m�x}dL��0׌Eز��j�3�B���B%KL���:��~Qtȵ'��!�s���͓u�^�VXj�LR�mc�5̘mq�i|0�<�ܤ���γ����%*��nn� I_��Q����/�"
��]]���2Ҩ�{t�/����wY]�W�7�4D�̵���>ū:���4�KO����yVDp��g��~��GwV���Y����B�6jR���16ʑ�8�'�+٠5̛�Io�j{����G����oe�We�Z]fh$B5��V>���=�<\c9��=�9R�j��P�r��3���Ӳ��V`N-H��<I�>�cc��s��\[OO�C����\C�((ʐ9�jU��V�d�|5����V �զ��C�r�Ms�hh>�Ư�P���`�	�������͙HŔ���������C����x㙄1�*��� NK��)ހ.���γH��p�X��w繒t,�{�H8�SOaH��C&�;�:*ǆ �5\�a�
Ծ�"�?\��r�E�������2�	����A�����h�w�f�/�,��4�����T�g�l� F'8���H~kc�sQ|�
x�˻�b�ҏFz="x^��ܢ�Vr�T�'�Q@�Y�����$�N�!���O�?��<�N��a�C��	����D�*k?����y?�L(� ]�$[]z�#��O3���"�ص�L� �P���VK�����\��N{���S�%�{����:�N Ϝ1�3~
i6s0Wy%{��Oa�	j}Q-i��G�|;O/�ש@�C�3��.X��WW�=�n��o�w�7ғm�p�C[���̸�ׂ�?�*�m���_�P4x%5��A���	�V/S��R�D&��dH�G�V_¡׉��Տ���2$��dp��X6����O�۲��{�#���� �r�����S9Px�BJU�L~���6��3H
@�^��k�����#x�ϑi���7�&�}3�����d�\e�da2����~A����>w��z��o:c^�J;��}��G_	�~�	����w1��
�:p���R����uDt2��=���c����@�6�Ѣ���|��;k��t^���� ŷR�.:+اO6��>�@�^�����CLm�soè�P|'��W��B�>��^�^k%V���8��J����V��<�ң�>e�+G��j�-���}�Cs��L1!���(yjZ���
RPC�T�}w��:���r�uv(�"��5p"ͰA(\K�D�Hnʩ_(�BxG�C��B�I�����1�x���"S.�܅��g%ߙ��qN���l�j|d	��?1�
�O
2&� P44��<���5_$�Ir�"_xb��YTH`�zX��=��G���&\x����O�M�j	�ug�I��xʟ[A����%�3��Oz�
�霜�9[sj�z��2��mqa5<`�l|��f��d����]ؾ������>�!��g[f��	Z@ڿt�N�w.�g�����g��rj,����;�uF��)��Y"e�.0]M���m����e�p��\)�ެ&a��������ՂZ]]��W��^�ËA`)SD�9��,�/���.��`Z��3��T�����b�Km��M���Y�.�ϛ�:�\Tp�o=��[Ծ'Xe/��տգ�Ȥ L�YM���4�!�dr�����ظ�@$1����ܡ��x	^�_��I%�@�K/��Y^��Ъ��	�*��nW�� 7af8�����Z������)�*�u�`����@��N;���� g�'��f"�˪��3�		�"�4@�7g"Z̕�"�����T��m�ڛ�ǅ!!�}���v䆾�ha��
'��B��㶔���򣔲4eʡ3�}�U���00$�}�fZM��mo@����~
�^v![��O;$~i�2��y���jx�}Q5�W��ub�5s
/ǅ�ZLĥZ�����"�ƭ�|��o��y�����k����t�t��9 �pe�B��V���K5.��ې�Y��"�d/���p��䉩��2�DQR�Q鐘��i)W�9��[��2~��Roso�2M�)�Nx�!.s�ox,�����ֵD�9+��,�z�XA�l>����V#�Q��>x!��z�����ָ�9����2����]��Fr�5� b6�Lu!-3�;c85Z��\yK:���
M]�k_�i|��w��p~밃H�l][|.%fP�mJ���0o���O,�;<Ed�����g�:p$�`l���`�̄�Z�+��d;�N���Dtg"�!z���"������`y�O��wC�f���2�?+����j���I�<�Q8�� 7�끗�^���[���v[��Jz�+^/0���a}-���w������K<sB�h%E홯U��6ό��*���}W���S�{m�
��/>��n�X���d��t�mm�>M��������x��2�b�b~���7�u���`"�9���o�{D"����J�י�c��{�+�d���	c��?�P�-��0/�1%۪��?��T(�m�X�/�D� �	�=X��-��]��8��1��_�P��u|R��a�����3� DՑF��e�c�ݕ��6��+�
;l���\�r�0(Fswe0Y�4��y۪{��H�h#��T��`�Z?ä��!oחu�*��iw� y+�fX'nɭ�Y�~F@����M�LH7=�x2u�/�U�W8u�	�od�]vK�`��L?�hJ���ѥ����-E��z�kp&F��x�d�>���)������zo�"4�Э^���a'D��/�#9{�{���>��n�˧b�vh��׹��*�{�w~���63�	n!w��j��^�_��+���C�&Rbf��%/��an���Ӓ�h�=ŗ1�̨I��
�L�y}��fh�ۙ�[h�ӭ�!qx;,m/�<�rj�^�~�� ��L~�����_���o�e~�����U53�h�м<Xy��GT��㮲��Qئ��A������*L�.�ܹ�?'���<!Cx7��D�������a�^�y#5o��>Y����󗺭�l�,H^���4�`��?��!P��U*��ُ�7��R~
��Z��:�Ĝ��<q9yR�|~ ��h�R�,�r��r~<(��ӿ��.��R?�>�.R��0/��Q?��n��e{��$�n@L?2s�qqӅO���_�ˋ�J����ǅ�8h���B;@�7�n2����$M��y;��|��x�88	QFy��-�D�23$b*fV�6e ���A�V����YG]S֭�m;�ķۍ���A��4��j��5 	��g9��d#��|��_�TğY��	(}TJ-�����O1K�!�X�F%�X�D��%�a����Kj`V��S������΁#���Sgd/�o���u����$	V�����)��A7�Sz���V����U_�!���D=��3 >P*L���lg��T[	��m�05��z�4%�l���ts��.��M��d
 �"�������lŘE7h$�T����j��I[|�wcB��4��qȇg�������!|�a�xo�"<n�dh��k�8�2�5kH�!�$r ����`'ĎK\�X�$C˘��9!ڿ�ʰd�c�DV�_����an�2h���M`'���^8�@��;D��ARHdQ�:0�O��s�/�M���n߅cw�\����)�Q�(��+��o�Z��c����7�[��.������Ba7��K"]4Pz���o�ufL�5g\l+}-��2l������#z�p>k�SO�r�t�gz�:,��h�~�	����o%�Z�Xk���]},=N
�ͽ�����	K����y}�� ��c�ً�p;��X����#X����X�7��a�r�� ����z�,�I맡����4?��O�b�pv\���oʞ�39&��0 >V�����O��G����bc��O@�H�m<1���{yCV�!��i�W����FB.KL�!v�W�����c�`�]F_��c�u�җg6rY�=�6�P�8�3}d����NO�����Z����
y�cn��?jt��������!Uele(�wI�WZ�č U���;!̪��8PY'���Q���sM��z�!6lezF���#@LX������gB��
��@|�Ü d��c>X�JlQi:Ug濪<Bƪ�V��k�����������0T7ĕ�gĝ0�/�!c�3~��g�/��^��>}����������>Ki���
���є�A.1�a�V��D�K=
��� �Y�Le�F_ao��=yK����A�?ٵ����b��O�7���
:���?:�%�8���6����_���2�	u���h*X�rC��E����j�T�PKw��)��"�@�4�Xr�$�?,�5�o4�@	�Ϙ0�=�j���t�7Zj�T4���F�?h.0�u<2H�zU�ł�e�Ҥ�H��,��6��K1��d��֞��D|@���9e�����Q> ���T���d~]����ӆ(�1/�˯��6^,�+C<"�)��*5�U�?�+��R�T�g�
{=1�X�$dB�R�sSÆF����
�˞r}�����]T�_�nm����9H�-\�7#lmG0Ys��PP�\��)Z�j�G��)$�����2#b��S$L��|�sxh��1��SQ�z�+�'o�$㗿Dk�ED��#�uyS��`=Rzn[�63�j` sH���H�|�g�{���d&�tW�_�F�ai��&�b9��}�eat~��]��Rd�@yhlˍ�ݠ{�P��������jژ4Q���G�-��-b*�)W������B�_2Y�(6@���?�hxa�����F��d��������㲠 ���h~}��rJ��L/����?��yZ��+�����t�w�/1[�Vh4�^_C�D�ɫ՟����q_ɐ=�5��0UP���!34�5ɉ;�Kd���W,�C=�Kx�G��:�$��ڑ������ɋ���M�����uq�U������w�Ptz�ˤ"�F��h$�J8&��\W��b�;�z�f�G� Zϫ���ڐ�VxӯFf�q�c��(�J������]���'x�E�{{�o^X�h
�����}b��Pq������!�s$?�q��v�K��r�N2�P��Yϻ�����8���^�!�֭�?�"�F�k���{�¸gl>Ifq vz��XL�~ٸh���ĝ&ц��W���2Vٷ��f��;��<WsZl�z-"o���0K�vi���;�P�e�~�%�O,�I���T��]H�p(��'��4%��K�4k,,�:�ͷ-1�45oB0�3���(��e������ub׸�8���'ޣҴ���"A��n��'"\��P3��g��K�5 ��x�#Ʃ��r%�Ѱ�ڽh�r�k����r}-��H_��E�
���a[SZ����3�<7�7���9Z�T�l�ִR�V��)yD
��IWb�`c������௚=��ߴm���+p��."W�Tyq�7��
%~i�� U� �fnX��/r)O�j�K&NT����#w�i/ܵg�/3
���H��=�w��͝����s�kG����������w���(��`3���>Zk��X�x�P�峨��Iy1 ����x�j�{ ����#�SLB�f�1KPE�u{n�W�JL�x��ϛT@����n#ק�?)fM�����[t*�W꫙ndҾ�	��
�i�M.�j���������?����o�) �E'my<�v���R$Fť'YV]�}ia|m'����QpΰYR\�W�>U1��4����]3�j�`�wz�/��^������%���=r������Ԕ��BA�B"T�,�Ʀ_�A��ᡕ��C��ފ�Bqb5-T!(L��N��v�.��pi5�f�ŊQ�Z0G5��Jٺt��
o�&3�5܌ Q�`��Sewu�xS�KR�t�LɥS��G�b��䬐��&d`*2	G�mR��yV-��!%��:Ts�o�����w��H�!���5��0�ӷ����5�M�a�vipP�t��	_�G=�\�d0�00n��-�ce����3�]T�5�P�K;�z�Oz��+�'}c�+�\���D�3�KS��9<@7r�1˅I���&YFM㜳��*����Osy�"�*D���:�d�@���]X���kJ�`��k�"������]��{��5;��/�D�5%Ҷ�1&�;ȹ�p�~��P5w��lM��G�K$�J���5�ڮ�����-X���4��+�h��WƖ�g�ENh�΢��8{f(�g>ˬ���*�po_�X���K�+�������K��_BF�U���k $�E�[�㵙���y��W�iT��h��hn]��9���%A�(i9wR�D��.��7�����p�Ke)L��W"��'���za�5��)!���qt�r�m�y�KW3}r�14�s؀E�4�x�2���\���E�>`�̼�i�{��p5W
J<�QoLy���� ���&aL�"U����苏��t��<�6�[�\9�CG������-T��$��=�e���>}�gz{����u�
�㔣Νӕ��7v$�*ok�aXg~�t1�\��HA�q�Ԃү�ng�.@�m;/��΋��I�%��c�
G�M�ǶS�'B|�u�ۤ�G e���&�5�a��o�MC�n��7_�Ķ�C��M�)���M����V��MA�׼z�;;�Y��%��k�k�7Uӏz.?�Dc%b���E(��8�s����ʞ7`qPR&���'u����o��/Yvr���h�|&��wz�|�R?�t����ڻϫ��2��p�N\��_�i�Ìl� ��]�+�Mي�B����l�d�X�m��-�����Z�}��|�ߨOU��eO�$�:
���w���'i�"[3�{���?��6��6Ru݊��>�``�j��1���	C�ո;>��
"pF��̞���/�)��Nw������8�����)����q`���;ɴ֏�Ȗ��Ƹr$�`���븏���E����<�)p�в2��X�u�'S}>��D@�Ō@���1��o�8��Ļ��ip5D	�k$��o�5��#��2ʆiB��	§�G�� ����:���Y��L[��h4��g�`yq����oJZ-�T5�����K>N8U�8�c��v�@��֭ �x�H�����k2!�G[��OEB��'BLhM*�ܧ..��wz���9�Ǩ�?O�f�k�U��Vz�#�������1�W�ޟp�Ϭ�xӺ�.�_���j����φR���o��XN���F�Q��kh�sxh
��$��/�R�ј�e��q��H�+��11��{E�j	�U�*��hG������vؠ��n��!Xd���dD�N�9�_%;jĺ���U�|�QU�����&2o��k�#��v�����B"��~��Y"�c�=_�_0V�Iy�;di�$I&�1�_8*BԿ�v���U�c9[��ʲ�=��q$�e��
�i�`p�zs���X��btS={��xǟB�F��9*nur�GT�Ķ�p]��̼In��|f��V�u�V��k�6��M�� �ӷ	4ǖ}�E�Do�+�V�2^�ӳ<�w����3S4�
��{]�����<@̅��}�d��0dk�4�8����Ni�B��Q81����%*7>�v�p�5�a cg�y�r�$A����Z����:5_���E
өq��b_U����e?����,��[��8�$@9��Jwo�/�`�J����G�����A;�ʁL��ԋ�NI5����x��娬������rJ|�K�9���)�֗��l�%��+[R�	�G���D�F�lC[��5��v	v��r&�&;����JR�*�\}*�`@����\�/a:��Y$dT꿠�l��Э�9�!*����i�:��R:uH�:�WDD{�Q#��]�%\-z�!�zV�j5/>.�}��mS;��.}�
7� x��Ҏ��vW<[���I�qU/1%�������)8�Dn�eO�ES6���zm�sw��Ur���A�Qgi I�����UK&�Ź�o��)�T\�h�_ ǩD��ej������`s*`����ޮ���s"Ť�����]��=���j���xMFC��S3J��d�E�&��0�r���粲h��=�L8���.���RŮ�~����� G'�ZAO`\���.�d/����0���Kӽ�j�F�����b�>,�����G���G.�;§��$�`���d"�ÓH�n4}�G�>����<	�0�1� ���"][����#�������aW�&M쓒���hʂ�/�x�/E�����H-y�o�d�S
��%�v#PX֟��5��?�v�#�88�ێ��(�u:og�|�p�Hɓv���C%���Ybǻ�,t9R?,�;j��Bٕ���.)�G�0s���c�H�@����Dz�!ŗ�
�%!T�c��܇�}��7�ʜ�M$�@Gi�?Y^�N�1�΅T��*��5|qD#�'��&+& �@@�m��Ndm
�\C�;~)t��Ժ��j���v�}�4�p�Kx,_��mzk%!=�g��8����` ��-�s	B���0�oP������������T
0[f Pp�)�v��hɁ=`�h�:iI�]흜���,�?�-$�K�7�.�qH� Z����]$�~�c6.q��䛾���g0�U8��O�?R'v�{u?�X����>���D�0TvJ<���}�7�Y�T�%�8�/ ��|Ҿ���48��snŢ��P30��}��P�r�(�+��<�Sw[<�*.��7ۭvA�KF)�tkŸ�0	�l�M���5	^�k���l���-����b������i�'{���/h�/f�>�
��+�^���
$W����ʂv괽��%/Za=Ƌ��=�1�尠��kQ	'��ᵆE��
T��Dh�T�	��bP��C�����e��|6�Pfm��¥f�d���W����2��|���;}�]	M^e2��0O�t>����'ln0�ۋ	��ݮ!y�~w�����հ�w�^"-�!/jl��w����rr0W蘮xs��k��#୿�n7�)��V���Q�VUv65�6�e���+�]Q+��G���J��L��	����h.��ǻ��@�^^�\�����\Vt��s�]����j��uw�$8��@�.O�I��@�[c�U��9YZM۹�(�E�4SC�Ji�hz0�����Z�����$�YC�p�(o�}�'���1�K
ǚ����W���GfIͥ��[0&Ux����m�XS[���Kΐ�����ޞ�~@�I��Ց�c�G�5Ȣ��=P������}{�/Ĺ��;���G_���B�����p�۪ڜ#���*���|����5�6?��h�F]��5�F���Z$���zXw"��^~ſ�a$9:�!&����qD�kx))� ��|',s�hw�S!���<M_ 1�}&����X�Q��P���I'~��8�jJq�g(����wW�APwvq}�M�QU� �*�0�!xM��F��F���߮��	�u�p�g�!<�����&QT3�(7r�K� ˏ��8��{���8JM��r��_6�#��W:�w�ޚ����p�����}9=��r�mėqC ��2����������Pl�á`E���3�K�+}e�E&��!�Ê�l�*d8�Jȓޘ�ĳ����9z��{�����ǜ-�Z��~N��{ҎY������{�6"�7�L�\���>G�k����(�d�Z}�L�n=��&�V����oW~���j'�d�ʳz�Y_h7r��ͥC0�.�B�\�}�L�y��""��0Τ���� D����(�
ҵ���
��/=jc���)P0��e�_"�>������:b!��1�#���:(Ȳf�x0oO^7���d�A�TLJ���MH�S9�>��V�a��[ �@�O�.'b��5��d����NH�1�"�X�%����2����' Ύ�� �q("����i��gM�����Ac!���xW�3�NJ-K��(������;U<ctm*�A_�Iʺ�j�_���Z��m�zCܯJQ��R>﻽:�wŃ'vW[�U�F�f��t�2pl�ۭ0OڿWxra�����������3@���>�������c�g|�]^��^�>\�,����!þѼ���X��LA���@2���2��
���5��ue��Q)q}���ƥ�]5�L��/���K�	�N�Γ���D�,p�p�o�a1�B��V�g'6gƅ�v�>��&b]�f·+�ub��o�s��2�m����@(*9�}�[b37�<��Q�*(SX���U	�L(����k�ҹ�����1Kr�`Smp� �I]ܚ� �$+��|g�L7Ϧ�O�} �8�L'��z:�>F&w"#�>K���a6�2�/׵f�����rA����>Rwfg8�@��oNS���Q����C�>Meh3�x��L�s\"��B��(Z�ie�%���=�A�ȀJo���`}�\��[���||<�$ϟV�"f�r���M2�&kV���2� ��aY���Ca��H�[e�%��<z����7��`^��(=�s��]o�{�S^e���_��*���^5P�JLx(�V���iX"�m�#�<�B�SPɩ��M`t��9ps����J|�4��pW�{{��(���p����wݶg����Z�H����H`�/���b<�:mR�ʈ.Pc��f���i�UVm�*6��ܟ���T����*�86x*'�m�z]zc�'ߚv���U=UD,�6�6�.��	�<�<�=/����YN)ǳ(lV~�B�A�=��W�WJ�tM�V+�qD�M]ln�˙����F$��S>-�M+dl�[H�b1߃va;L!�[ٵJe���U��:�&�G�5c�h^ê=M���0�Fn���.Ipk���g��xK�3�0w/sCa�/o���Y��2�-�t�L�v�?	�~N�i�g����:n�(N$Hc𸐁�0��� w����®��	�{Ct��� :��H.������R����AŲ(�8[�k%���~Jؕߚj��酐��j7�4V��
 sUi�(jy�(�!>uⴼr�>����KD�D��%VV���[	U�ӌ�S�Ì'�M����N,��>���q]���|����$�F֮ymV�j��m��gP�&�������(<�̳)����
#s�B`6�=��on}�?Ԣ���[� *p�_vH;\���#7��u��K�z�I ِ�2\5q~~���i�a��G��v�� u�ʫ��
��e�Ѽ���G��k�\㴧_�.��zd���G��]gs<ł��:���J��ܤ[�1����yBP57�k-���4S/�w�t�\�+F��1�$��j⣄�$U
".7Ev{���ˏv6灯��X�
W��g;��m�vuܣ��J��?��/���z���?�w�41�f�#ry �����mlv�����ߜ���U/�L�8j��)JN0�O��������D���������Kd�V���B��y�� �D�(}Ղj�mra�:]-˃�~��;��:�u_���p��4��&�.y�>�/�]��E<8�6')��eoBs7��׎WL������Q�Q�l��Κ��m9��	��v�u⅍{M�Mi��.ߦ1m��m��ʻ΃�_���R�o�6XC�q���o��mF˨�+��AՃ�����2}��@�[:8�V��k� ���Q~d��	S�C��G�e,�y�%�D�"���<`F�+w��^T�}����@	���L��ͯ�~<^Eɠ&;�љ�o�9QJ5�߂�.-]�^4\<�֦�u��L�Z��x@^B"�%����� q�kλYqV�Z[��d$�BCN�9�����Z�J�Æ��T�,n�t��"H�:䴉LsэL��n�ȵr(��n���,[�������f鐍��%�dY	����ކƁ�@��aN1u�+�c!2���=�1OC�-3����9\�eꊎ�5��B˞���[��if�O5C�+/l7�P��HeX4��M�t��=;���԰�'��T_��Ь�e �I�2a4��~ ��2e�E�MY�D�����aW��.j���r�������I+T�HcA�k	@������gJ� �Q
�V�A�9ܙc��W�#��
F��h~���ƶ�@�Nhy���h}� O'T���|ؑ/F,��i�(z��Q���$=� �.
��:k��b����AmBxf�o[-\�m����eJ�.O�/#O�ζ��-q�r����e=J�8��̀2p۲PJ�kP���ӑ��/�.�K�Z�xY�C�q��f��w4�.�z�ή���E�����Zj�F22+���$]�����ݙ IPtn��̚Y��q�tlE�Ìj��9�K���,@ϛ��o���J�/��z�A�:I1��B��O�s4����K�	�U�=%_�4(�֤���]��?[������-N|�|��4��yBkzL5��[��`�B����=ѫ;�_	��+���<�%����D��EB��0���"18O�i��X��FtDM��ˊ��C�w�O$T���V��瑱�}�6�gq���A�y����TR�i��4����<�[ 	,�p�_
�Ï�<I���^94�+�W���Ζ�z�'�����O�M��,��_ST�ŬweG��i�Œ����X-��f�U�������K�j�qe�F��]���v4������W���InBT�����
�/_V�������n~�nsn�N��f���"��g3� �t��O��T�p%#��'��p,�z�uX���[�Mzwڛ4zH�$���E��m�b�v�Ru�X�'�cI�'��)Ry��}٫K]�=  �,��m0s�>W����r�4����a����Y8�P@�>���g^��+�4Â���[l��B�`����ٌ2W4J�6�) ��4SB9���{����A((��W�]l9�y^��x7�P��W�2�P����(��n��tNXMР$��믤	=����F�f�c���]@�q�(�$��Y}p���C���~�s�n�`�g^�%0̐��h��s�M1N��$���W�����!���3�5t�����(�4�2�b*��ҹ7J���p*����f�u~�'2֫&�="hJ��U,�y6;K"	��wvŔ���Y�#z�%QL$�2
���9�;J��t��6�ߤ��ƋF��������]$\���Z��PNT�p�� ��K�W���TN���6U�ީ1�)��2l$�� �	�|Z��D�!�@�K���\�eY��L7������J����������R���#�P����X�}���5U2�4&榶z�q�t{K�4{�X?��ճF�,s�j��<�Z:nJ�~���R�3i�ˬ(���He֚�.<{��wܠ���!���J5M.�h/�����F_��@��Q����U@��2(��EsMW_9#�ו�+�6��v�s )�؏���$��w]"T��˼iR�~���V-C��|[mӶr��Z1�EV��
��>�p �Y����Y$�_���ږL�m3����{?J;��"�_4�@�$�i>!���B�,uwo=�릀.P��4:w��.���_|ؖO�9ߥ���
�R������(KHo�ڢd?kJ����J�n�l�7k@#ш�-�gx5��p��T$~tV���ԏ�X�Y�UJH��׫��;�߸ϸWPyGk��b(�ñ�s�U��;�?(N�
��2~� ��b+�r�7�I6���]
�;>��_T�eɒ�'7�O`�bfpқ4e4��^�B|}�N��L�>�|b@T|�|�|����Vu5-I�AZ*`z�J��/|��]���s� s�{���s��#m��O	�E�W�o���jaB3����<��ޜ*�1*�8��S���b��ߧ[�P*L�C�_���������z]1���r<�h���
�����qL�Ѥ9:���"��+剼]�J۾瞶����)w�MH���S��|Q�a�*U�`���0"]�eq��c�i�)����zIR��UH���&���Rw˱��WTP�]�~e�ق[*#�
\6�Rfn��#�n��&�#o�o�#b�S��X���Q2��i- M;r��j�O��,1�a<y��KF�+�d��Qi��ܫKkOy�$S��s!�����I�ί �,��Cs�v�獫0l�rr��A_��/H����;�[����D���"W �����,W�T����k�i��8������Y˅�.L��i[_�֟ɋ����|�(�hSa�괍�9��y���#�{P����+=鴼��4��Ys��h��JE�e�x�5�T�v�V}�2k�����{mE�ߩ�4B1��-v>a�3����
��:�:�mb�υZrb=/r������L�ݓe��;��T����������?6ō��Ú��4ؗdki[>Rn��'T�O�$�v������/!�rI��E�4&��FF���K�m�琡�Ǣ�>��&(L�p��Bç"�s�#�b�� �X�R�?wW�.>�\}�b�_Q�K���g�C�f�G�X�cb�.�a��rG9 ��=R���� ��#fPr,���v�v����m
x>��٢$����#!��urSH�bF�T`���V��8�o+h-ČP����O����-�q�D��J��X�Z��¬,�6�B����&L_����sN%���D,��X'��HHe���Sh�(4�� i����G�>���-�`�OYfA�U;ն���
D�3�����hK����	\�n��Z`�4=�^�;xx�w*l����]g,�s }H �w t��f,��#I(H��Ú�g�B�j]���E�X¾�!ո�G#�x����I�y���I#��������6fݓ�_k���6�h~J�40o����Km�T��!kw�.yjl>} 6��G������O�rT�@����[[��|ѡ����6�P�5f�yZ`�Q�e4��,v<��3���N �M*�M�o痴�)eC�Q�[J�C\ץ̕,!����G&����(��r�^Mux�n����Omg�,d�ד��'��vJ�����:6.��ܤ����k?�w½���E��m�Y� �!�5Xг�F�@��֨<4��u�$붦��!�/�0��}�`1P��f7Q�//V���ང~�N�,9i�������\s������j~V�s��Ȃ�D�~�{P��lk���z\��LNN�g4h�)��7+KK�� ��q���{=Ip�bq����-W]�O7�vn�u�ќ�r��G���Wx�i���#c� �صZ�]䍱P�uUUlUo���v�n��i��nWԤm%W�x�tv��C>Y�k)�!���G�"	&�[��(9���Pwų�R_a�d�]�����g���7+s�w���3�)�Gnr��� ���;�v��1����/�9!�ι$�[����]V�#\��[����\'u������?��8�|6���x�҅n/w�5���i:�\f�Ǜ��_�M�5�n�Ŷ�O�>�CG}�aF�6|�L��';�X��.��'H��~U��F�d�P���Y��u*�#lF�}��<\'�֯����o W�Iz����$7��9�/:S	0i|�քfgVq`�h�"�
0g,9S�>��=J�
��'���gW�y/�WR��������q��w@�����E��������y\�3T1�U,��~_���"҄���'�x?�C��H�2j�!��Wwi�4�����ķ	ғ�r�����A9V�|ն��f�#���&(PP�>S~D�J.n�8�&���e�v�d1"���B�%�zq��D	�u<�P�[uΘ;r���+�e܃���T��`�=�_P�����l�B���3��N������xҁ�b�w�y������������u>*s�yϜ1b���=�������t)��p0�J(�W��byMPu���XJ�g��es����;��Ǝql�~� ���@$Q�|!p�NM�d}l?�h�Lu���_S�7��AA���Z��1��	d �MR_@�Έdă�5`��3.�1��9�sFdQ7�og�2"1a3�X=(���WZ��]S��W�i�>I��M���.r�ŷ��4`{s2c�T�q;���^)]>���/БZ�_���k�Z�_��;n�<��f���VMM�yhɀ���=�IiWp����A�P�
?���tQ��ɔ��֑�/98Q��jzV)�Q��7���!�yL��D>V/ݦ?���$p)�=XV��hg`5E�:X����Bl�E$�����58�z�kn��q�.<#�_L�O]�����7]�P��\:�H��S�*`O���|0��Rdu�~xG�GFEb��P�$6�<���������B� ��jw����]�j�X��UmuF��|l}Ձs�R��һ��z�0���X�0տ�͘k+�K5Rԙ�QiqY�R�IcG���v�h�s4��޹�=�|�}�\���	Ny�K�����<N#�}��5�����h�ӏ��=twf:�_5��7ut+s�D��]�I�E�Ӛ�]�E1X[�pC,�"bȤN���jo��v�G:\h"����? Kܽ�.W62��o���ѳ־D�\q5E��x�x{5c��k�
�L��;+���9������ݗE%��]��"�CX~�x11<G [i4��wYme'�L�
��:����ᠿ�A]��X�� ���^��!�b�`��C�o|ru4��z���< $�_��xPIg	7��x,���3:���)5#`������^�O�TRZJ#�̉h��j��
*�aS�e���y�Mތy�_�\�y��+�!v
۸�:�f�x�"���p�f�mUV(�FkGy����!ߴ�Z��*�����X��iJn��y�����V�����#V"�@�#�e1�3����������w��0���
�d��4����@5���w_T�Q��d;�-����:�|��Գ�����4;�5�kY�+6���R]ZX�NX�X_]���ښH�A|���Y�#9DO��I�N��J����X�#^Z0+�_�=�R��[�n��O�]�������� "��Zo>���9��^>���N�B+2¯�i�l�܅(��W�4���g9��0�]L��Ј�+U����+-|��asu��8�G�[���XUz�t�C�����oԗR��sJ^x<�3� �W̷��Բ�T�.��.~ �9�٫�uQ8�f���)_dS�]9qt(�[	��V]��5�{��-������9�^u��3�7�e���rJ$��%�8L_���;����������.��F=l,"j3�ۛ{� �n�,�a�A�Y��)�x��s��r1�G�t&�e1�wt�2֢�0�9 �B��z�:�H"���	��}9�(༆��@�y��B��:椣�$s{#�G�&J(<o4Y��U��6R�0k����_h9��d)���{�tJ¹N4����0W�I�U�)�4�<h
�����nI��h���N����qٍ������H�B�n��+`;|�����ߏ]h%�x�Q�4�Ja
��-�@�,u͙�+��Qӱ"f��v��1}��">U�W9/ �B̒r�H��?ɍ{��B�.�֟O��(WM�����F��}��`�fåVس�V�f+w�ՇƳ�1�-�`w�����)�rUV?Mt+6�Z���6̅��]d^��aS�~��i�J�I�A=.���|��J�o���J�Ռ&!�����D�vL��mSm[���׺��Yﵓ��V�&�4���O�.�����n8�(5��0�6ĲJ�I�
d6�|�9�!j+rCt�r��zS��M�}2�
қteCO�x<���A����o��-�;�u��g8�!#��/��
�l]���6�Di��YY*�*�5`83��B��gw!?w�wCX탸k��� !{�#�~���������x;[�|SS�f���н-�t��(����-_D���]�>0���$���*���Ә�"���4F��zdpUNI��P��4�pL��d4ү�[W	����K?Su�'�Ҫ!�Dx�����)8����B���DW���=�X���O�[���-�	ʏ���+W�b�4��G�# ύ���$d_c��ԋ
��n��?��9�TXj�G���#�)��4s�����Zhv��K���ԑ �C��
r�̔<U��;�|j~� ͆���>D%<�_7��PW�(�޵z�$������6�0c�V��bż��[ie�	��{w®�MR�T6k*��mA<���`u��P~#M��b��}U7���I�@����[������#c0Z]47�d)�~��ʩ��9#��?>u��*�%>�:�cK(&�]݇��xRy�h��x��d+�י
ލ/�,*�c��>��h�F�`vɈ#n^�&MVL�����<O��4�*0q�������J��t^�J�3�@:v�����h4���Vtk�S�0�n��<�"�"�sR����E��iG?�e��׬��]�~a�R�+�!�T���y?�<���MzBLQ��:�&�)Q�*2fIl�{O8�*B5��jo�� m���b\vR�-]�����n�Y���������8�W��u舊ixyq��Ř��S [ZfY�]�JI8ʥ ��$�Wp��.<��(��;���˝��ĥ��5�Č�7���.����l]%�?����� 0��,����t�o��`6)�����J�$�_��2��B"ɧJ2�G�a�#�����YO~�I�nk�t䲖:���PY)(��.aϛ��hj�qd0 Uq(�9u�Gb�Q�,5U�������iުc(�����Cſ:�E:7@�	��(+ -BR�q�BU:Odg��[G�C�^zL>���fu�ByҞ:{�@�{�.��m�q�jwI���1g�Dʒ��ÒZh�J�.�����4f,�#O����A��avz�a(�4�=J�R�n�I#��.ޡeNQ�C���qE�w�Z���peׅ$�]� ���V�� 0���TS�񟎎><���}[|Gp��9�k��D��L��J�A��G�<9��Rܓ�4f��רM�>��Kq��J��ߺ>x�
r�6�E坤�o*�C��6V�i��A���k1��{Ϫ��it��=أT�������ʷg����/��.�-=���B��l�ٱ6���,td��&y�L��FS��Ukm��nXΔ�lb�'�V9m��Sn:�m��X�4�:��oɮ�� �B�<�=n�qHyU���F��p��P�W`D��ѥ��M��q�ŵ3�h2����s��qF�\��a�m�tkW!T�4�x�3��'��[�;�^���u�T��Zcec9l���Nܒ��;���p�S����βi���R�/�#�9��sDq�*W�O�ǟ��\N�ʚ��e�h	�;ĕʶ[��m�8kzb���+J�!)o�!�Н�l4}�|�l��e [���BJ \?�?��۟�g��Lݬ4�����O�^��33���b��p~�uh�8� 8.e*�*��o]���x����52Z@F���U�[^��|�V}�4c�(��p-&�Vav�@�'k�~t����*�X6��\�-N�<�_��bf>�M�gq������q��:�_n�8�%��cpg��#GR��d@Uk��7�A@�Fy����G/__�{�J�5�"��:r�u�ќ"(�q�tē�.��_��#�m�l�֓�zq'�d2�7y�j��\�#EiC�C�y.�3+;�r�i2���Q�)�*.��g����c�кGɌ�X�����[	��6'��8 �шF�%���͞�a������F�ý�X���p\�
9�e�&Oy�s�aR
��4�������[:#�Id:z��~��Rq�C?)6�o�݁u�S�bĕ�<1-�wz��-ZA^c�A�N렻wjH�L8�Y�Ы�R��D�U:����F��*����M!t��+k"�|N�l�bM�X	��)��,���ZO8�Tg���*Z�2��S�2eÛ�A�^Ļ�l�1~f�QW0���z�źd�i2Kgo��TĄGņHƕ��*�e�?`�&F��Qm(8�*7TP��=��7��@�揍nW��xp�*��d��D��'�Ƅ@����Z�?�b*�/�=~	ħ��I�Zz�9�%^�ꂰ�n��pk��g�.^֗�B%n7ɻ�����}+�&��
/�R�x�q�5s�C�g�EH���z���� � g63қeɌ-sx��NHS�Ix�9�Q������Ϸ��8Dm��qFR��xy3��ڧ�&�c��aZkɳ����y��s10�3vl�(�mF7|L�5�$n���_߭�)3.
扳E#U?�z �	a������� y��i*!д�(�&�
c�a��&2��
��$�VI�}�C��{�<8�z�dL{��+`���s����ǡ9d���eL�����،��N����X,�hߡ� ��'�t����>������v��#�K�PX%73�ɂ���׹i��������=�L5���?���okQ?�z�Pu��h���	��&�Ay���5Ө�{�8����#���1��0`g/�*���VfvE:+�3�5]=7?S���#Uo��ׇf*~�ʣٌ膌(Wx>*Κ�QC��r!v�}8��ECV�ӈꄡY�	i������g�H�1��@�[�4Z�Aj�����h��iӺ�,���ps�Z��t^�q�I�8@��Cg������Cμ��m��l:�:k�xxt�� oէ.3#��@{�y@����%'�2�Wu~ga��l��ǡ86�Ў�.��������/���<�_��]��(���6E��kuW��,�c`>�jW��Fs�6���^]X�
��k�L��w	C��dF���4/���#c�>�=����q���U��Ҍ�G̿9�96Hsc��V�����4O7�z�4a7���0.I4w��K^�uB���r�V~��E�y�"��ZP�D�y#���0GWؒ�Z$������ 
�L��y����;C��z�:�2�:�=A�Ǣ��9�m�Ϙ,X&���BM�I����[�'�ط� Q��=�z%aa
~2j]o�>��G���I���j�WjXl$�u2�-���@E�j1t��t���B�9���ֱ�~*�=:���y�	j��l�*�����hb7�7�B�}àOW7����38�k[��\�m'�=�m��$�0�����1?�h_�D'C��)�?�.�:��Xx+�Ԟ�6����9��!���Rp�1�=���2yc���x�O,�2p#<H%H�r�@������K� �2..�P�F��|n��H=Wu�ag��Œ�gq�2n�W���-&>8@_"�>�-�DY#W!����*y���f�����:ǁ�B�_����=��8��KU�h�8�FP!�s1�DeA<&u�V�s�p�"���@��6��tNL�pQv)��V�H���^�9\�7IJ���J=�k�
���dD.��U~���b�O�����J2[*W�<`GItM~}?�7��h��w�7v��0.j�T�DS58n����eN���9�t�~
1�6��R@՚{�e��\�pjg���hj�� Ӝ���"��\�WGY�ښ����2"{��ėg��E��#E��t���/X?�ρ�Ulh�B�9[�qΩw�r�B>z�I_�sx�]b*�����~�/I������z��jw7�U��3,�NT����κ�o�ظa� k;�K���_�;1\w�g�pZ�\�+��& �#�g��qT�km(v���p=��|�����m1����O�]	�o"��=@.���'�l�G���Y��o!GP��㽏Cg-���،��]L*o�v��c���sc��˷��'�X�EU.[h��J�Fz��H��ͬ���DI��琂���ʑ��G����9�=�I�Zߥ���a�ߙw����;�/��3�}�N@�ߏ|W%|6����h=��%��l�i��Rs$JB8aO0G�\xI���V�Cҕ^�CE���XRvvVp\j^u�`�s���!�����~��U7�9�L�iCoD�󞷇F��1'��"3�%���LyJă�"1 �8"Ua�3����G�'ry�њ�
ZD�������6uy���u��l~W�r߳�v��1[�}��L��4;���H����"/�zH���H~[���gHVF�i��'ۍ)�3�� U���?(����zU����wB�:8�9\R��Ν��}C���FG@���v�A��=���C~4��8�̑wX���ÓU�)'��ĳ�������o�@^���]����e4^i�`�5--^&g�x��
<����)�����p��|*Ȉ����p�tW�2��T)��1N�TIo���D�06W�eqd��É�(�;?u���j3����
��ׂ���z�#Uu��݆y�:�.Ē�u(U4������F	r������/D��<�Hں�C��RA5�yq3�=2J-��T�tʌt*r�K�dY�,'H����[�>&8�� k�n� �B�HƇ̿�?��R�z/��T��$z(��=�z�h��C�zB-��2�vO%nu�A�EI "��X��SBd}��be�-�\�m*�4��w�G�2����)mD� z4�<����L` }��{<7�/E�J}9d���=W���_\�?];�4��������P��W7^����8���"
�<̠�&k���"x\�[N��,?�c��>ڦ�l|"�z8�L	q'SgG�gؾ��/�Q��b�|C���v	ۓP�:h1�}~�Jvh!B�u�ʘŴ�K��;���zt�GW@B��H�H�Q`B۰�]N�
��hɛ0L+��5X�8��`��
�\��1��כ��{���:ma=���DG�ʈ{WU�߆p�7P9Y����} �f9��h�B�ĥ����;+�b�r+��0a���%D��������8�Z����NʈxX.Lڐ��Tf�&d��yY��Qh��l��Ev�]��*ƻ|&-�\q��g>�q.�bHH���������~w�ǹ;��p}9f��?S9K��g~7��f�ۯo�+͛�$KR(aY����57�];�����m���U>�d�!\�!���2� 8��w嬀!�O�����	c������"��c"���������^��t��y�8��I�	˞��F:O/�����t'�P�'C�/�ԕ�nmv$�������w�iJ}ƴe5�z�fI8�A�Q����ϸ&n~��I���J��^�|V�Bِ��]�D�3\qZ�cN�'�^T��m��9���)*-$/����3f�H.�&�d�G�$� +��g}-��[��n�.��L��Tk6�꭬�&B;�$J��'�P6�6gR���=UI����W��{m�Uj��׿G�v)(�=ORp�8�������yb+�����?����9�Q,�O3�����S�C��X����Y,2�h�)j�䔠�<Hǂ�>��i��Aq�̧ֱ�"4tն����dX�H7�}U E���1l=.�Hkm�j��-�b�eD�U(�p��Ό?Ӑ5�iR�>J��h8�����ی����b�Hr�+�I�b^"���j@P�[L�t�2P_bdq?<��%-� ��+���?ܛg��<��3.� ����li�˹b�N��#�3{��7�U2�N�b���'�k��bٗ�N*����(�g@ q�}H%�t(n���Y'�-ޑ��@��Bn���xk��2#�F%\14F��C�ł�c%��j��zՅϳb'MK���, $`����ZЦ�������g>,�wrX� ���*(hY�x�.�8�\ �����b�C�O`ސ��$Nms:�%����\�A*��6!�c�^��4?����~��@	�(��p���1����9�@��->��˓���tk����&G��c�|��~�˓�
v���>��8;�+����Q�i�������"��2��#+zd�_��+U�i#���+� �ʻ�)�$�w��^�@���o0���[��2E�4|j?A���tm#|J#K7���uRf����QxGJ�!(:�kc/)~�_8C	7G�8~ׅ�;�(��<Y� J�d���;�d-#U6�:94%Љ7J��C �j�R9�Y��d,k�f/��(&i�q�`��j�V�fp^��Ê0��&�)�t��W!"��ܖm����Z���U}����Z�]�v�	��~���%#���WUZ�){>&�|c$��6R��s����j�
H6�c��
��X�0�X1ˋ��t���n�	]�Pu�HJ��9��|`
�ric�^�lSi�V+`��{��#���V������[���*v�
rG����c�v�K��A#����'��ك؝(K��Z�P*�B�ۏ�ɸ���O���m`R�	�wdc�$J}@E��d���u_���i� ���7ۙ������e�� Ƹ�Z��0�x}�`Q竧NY��ÊZ=Υx;8A�J��OaE�N�͌��1t�N�us�{���C���GI`����3����8��췲5��q�oAw.�/È�L~c�-
�_�E
G9P,�⁻"(���&�h�ub�l%���S�2ᝧn��@�9y��;�Zi-�G���>���UFPmf?��)*Gܟ�~�`����-��)\Ȋ�5#�^��&-�;�Ee���M`��rٜ�ǘ�U��SN>���|^���E�M�,�Ng��G�m_��9�&<���i�G�A?C��R���K�ո��k:�^BL�+18�%ug/5a������z"��Y�m4X�N�,Kz#�d�,�
�dQmI����us�[��&�?h��ݸ@>���[��RjM�0����=d�S^w��]�V�2� )�U)�����Nب�*��	x������js��)���I�,�e@���Y�i9�$���7�J�D����+]����� ��&��j"�eׁ��T���j�^w�y�j��0�kԆ=�M�O8���Q���M�(�lFA�k�M�hXd�b�y0��-�͜OV�$�&�p=��`�^u���̄��.nwD����o9�������ѣeI�7���T1S_��^�,�+ȩ�t�Q8�.sa@�6���4�<]�	��c�ʇ�֗��7����>����T� £҈��H���ݶ��V�:M�NתG����xU	 t�ʻ�>c��Xgu��U z����ԾP�!�Iխ+��k~�`���O"Z�UNm�;�a����S��b����!h�*��9��FlhN�����{�� ��׀2�;VI�dN*�{ɗ�"y�3a�Te:8;J�"�m�f�{��Z�L} >����6_ȟ�f��
`If%# �!u��Z��P@�b%�,�fO�/A��9���MP�b�)R�����,;��Kȟ`�T�]� ��*�'���r�r'�H��Fx����]��ͣ1������7��4B������/g*��a�۫�L>J}��9N��>�-��g|��du#�MIIO��k��y��H�k����7;���g�LN(̲B����&�u�P�9����'�*���.=-X�)Vm-��K�^9�c�r��k�
��G�Dj!���8f�/�B�t�$y#�6�NC��&�.f�9<ua�˶mH�A\9|�V��2�]�Y����4b��Z�,��jtҞ+؀Sv2dr"mΚJ���2�J5� �ɹ�W�S"VY�����4�kl�p��mh�`�q/Z �e�F1��_q��s!綊O��E�σiK
��О���@�^�=�� �i�i��_���Ζ�Ym��K.CѓALG�WX�&H��R��_l?��^���=`-��{�oPRS[�}�齫S�;#��o��h����	P�M��!���_��[�f����r�|�4�_���gb�C��#8?+�o�^`%��� �D�9�3��%������f ��/,�M��<���=��@a�K݄G�9��0���a^�Xr�?��m>Qe6)��0=�Ŕ����y)>�cn�q�3L��ې�^��2�V[QF���Ե�V�+���%�D +� ��0�-&b��h�;�uB��|B?
�^ѡh6&C� ��ӑ��4ұv	�|4ekc��Um��^�WێP�l�>,�eB&���ܶM�I=�������j,�"���/����U�<c�ÞM(�(��I����e�2�o6
>yj�r����`��3)����j)�W!qac\�~3H��,r�ذ(l�K8�:��'�r�k:���o��M�ъ<�����X?���l.�ŏ�Xb>�bK�x>?+{�Y �r�fo�a�ZMԘ��i��1R��,-2�8Hȉ�k�|�*�	X?�����R�LY}P&T��9�ِV}6��a��[��;$�N��z�����q`~<W߀2���b��G�X�B���쬺b�m䄣$���݌U�mr���n�"P��\+��6Y�GSkyQ�#3�ͩ��9:ƾg��0��lyZm��✠��Q��@�u
���'ȞSӤՙ-��I� ���e�j��L 	�<�Ŵ2�y�5� 巄tN����>���d�\A5�_R%��G�C�{�;������f��?9qP����A���e�O��1y���y��]�~IU��E�h#ʉ�M������A�K�
��	�e��R�+RF�Lz��W�7���pK�R��9�~��+��}{^X�D�=�S�R�������1*2!|vC�x��H$"�,�u��#�6�q�[\m�]��s����<�f�>�W^�{�{�~V>{�O�����ɼ y7�Mطޢa�^R/)~��tv��B�^.2e�oQdJ~2H���T�����Җ�D<8Ш>ϰ��(�E:�~>�"_ ��;y$-�*?	X�W�yE�h@d�l7c�0m˘��'�rI����$�	�o:Rq�� сE��w��ѹ%�� N|2�%X�p(B 쏍�^��B�����/=��5��32�[������o�8y��3��#|�j�ۺ��m��6"��h4vkk��Sjf�%����)Q����C���c���_�mQX�\��j���0]U�/�NX,1BPlΞɧ�alG��[$���ޤ�g�>Bp�͜��1�;��N	L)s�7`I���P�~C:
�G@=�cu�[ce��ͭ��r���E'�q�ȝ32�6)ʚ�$�䣧}��|����;iA�j%2��0���[-�%�ŵ���]�C��b�A����' �F:�O�8; 1]l�".o�<��@�J��Sl�+}H�z�b��,G�~;-��Z�agLڣ����E�?�4�ԑ��5X���_�O��䰥��-90+d���<0M�2[E[�|5�B���n z�������΂��o��Aꃊ��I��Ngn$]�¦�N���� �5)ͨ��l�U9ƊvZ�<��t�%h��)�dF�_-�� 8�O����Xs /���c�_���;~@�P�'�=�c�mY�%�r��"�U<^9�|<!��"W�/�o'~t�IOy�0[o|���� ��?�S�E��+�����g"�:���N��y<`�H�N���p�w �>l���zI���M뚅�)N��|�����(�����M^|�q����>����%��֜����̱u�W{�h�;]�.Oׯȃ�v��#@˹���(����t�)����n(	*�lwmc�[ :u�9���7�Tfj�7�
�X���y���tf	�'ͧ
���?��'w#�Ku�R;���3f��Y���ɈVw��ȃ[��Ø�4Y$��|�a#~�Av���C��l�.d?�VaX�`A�!nq����j/����+���Y���9�9z�Y�l�8�Bx�Q�m���1쓥u܃OZ�*G臟�R��_	�g�.��6!qG�G�r�e`�uwo$�ʛ�ê 3��G>�����;|qY-ex�U�C�;Q=��|�w\��� a��:f�<�[�׹ǃ����r\$jt��v�/n��JF�5����5Ns��A�4,[�)fr��ABT~H�ry��FFZ��jS��c�N`Qr,jsO��g�ݛe��:8�R=�/%��9��ò\d��5��T�B�?�>����;ڟ��X�NB�v�M�����[7����|��HXV2[,��s9�}�]ɩ1�͓Q�&I�0d��y�CD�$f���ȶ�qS��������Rܒ�ďǺϠ�PHݴw�|j%CAP#�~0�\�߇�]/�i u�<��0=�s�����9]�k�c/��M�~{j��05��l��D�Ő��h��J�:qh߅TV�a:��p�7E(�Q�'�\�Oy���T���8��m�/�������H{���I0Q%L�'
���V�+��s��M��*���@\��#r��R�WEj<��?���ѫ�Az�8����9�-!�M�{A�O�a%��cY�G�Z�4��*a�1߈�{�<�Uy/�1tۭ�����j���M,ù
��z��n��;Бa��8тs��l�3�Q��Ιp���V�nb�)R�*~�����.L2O�

w>��_s�$d[�"�(��[��Q��,� }�:�*\9�����p��	� ����H��s �p� '@*��Z���X<#��L�`s�ve?炦�EE^r���y�p��aU�[�Dl�FE1P%���Bg�)y�&�s#O���u�W>,�*����24Ӳ���Q�\{鞬b�V��APKF���|�u��	��~��$���RNA�9�՗��]�R\5���K�ϥ����E�e��7���I�zr,�+��v@9��ڬ,��K�K*[Ip]�Z�=݆�B��M;tð%L�|'���������o���w[#bF���9�a�w<F�SSK�=-�`߼'��dwEH�&�֢����>մ��Ԗ���{�:�Z�f�2]Д~~��-��/1�e z���E�K���q%q���}�d��[}��Ql:��Ѭs����A:�����i,�D�@e�ѣ�撧���e޹~DO�J"8��]+��I���&g�=9��6��)FY.�ԮS����%,o��E[�K!Pd�@��=~�[7�5F�Xi 58$F����� ?�������l[�p�)��+���y���x�-8����t�P��*�1y״��߂�����G���\�\I���Ս�ɾ�K�*��0�MK"�{*n�D��Bj"D=��&�.hn�ֱ::\ǲP�b4rB,r
d��ܐ�:����_7E��+D��r�2���[�e�h��^��~rà���_��UoԤ�J�`�B%��Y9A؈��A��T^�Jj��cSkĆ��v�Ug@l`��y���Ե>n�����6�d�U$q���	"`* �P�J,^�uo��w';�XL��TK���w~
Ra�m���T�;vz"MNA��E����Z"b�n���u�Ʃ��+���K;9�(�؜�_��,��gC3G�\\sc�l��i�Ǝ����G�X ��'�\��~�/��eI�� ��>o�utx��u	6��S��<��՛s������>j$(��۸FqϦ�|{6�
�"�eM&	�%(_(ǋZ�x]�H���G�q,�^�ȬS#F����/��c�U���=�ͦb��;���������ٯ�:;�5O�\l|�UA���\Ҕ�kb��E��,�c�R����}����д�E���ӝ�q�a�#�Y�Cz���}�EV�6��������Z(�G�J_~�.�;ˬ��,ZM��\�JX*!�.�^��M��Mǲ���*������-Ŕ��
8!�y;Df�����b?af�P��xk���R����T%:m]2���%�����^';� Ń��^��+n��?9����D]���41�װ��G��8�p
��G�"\�.��P���XZ����f��jz3��F چ���oSB*}�K��DX�J�A:�:��K��uϨ��
/�O`N޸��sB��@�(� v[|Jaj�M����j9x*�`&��Nt���[�'������z	�����xTT?�r��Ϛq���uLw���&�!ą��B Fb×5�3WX�Hz�3�K$�����-ڟ���YT�Q�f�ݖɱ����_M�,s��Fy��FEH���T���X���#�_�5�C`������ z�uab�@/b�Iss(v����o�q�,>9�!�����Mxj)�B@�%�aj8���u��r�NP|r��p�kBF�����a�t��h���@�ϭgΣ�|X�3�����V���Ī��~b��h'�C�M�8��H�C�V����
�}���?�a��3�!�й����2j�']D�P���	\�,@�zMh=�	��)W~r��,���������Gb�0�+Y}1���q�V~ Y�vK$���5ɔ}?,�B���q��E���*T����o U(���1��m���Z���'�N���ۃ|�9��u�n���Ũ�X:O<��c~(�S�\_|7�U���]AX��UP��n�->���W9��m���x��z{� �;�`����Xd�4]�>���`��ݮ�F��)�'%)R��;����r̅0�zrs(�8|�������gXӳ�?�N[������)i��t�̻ؔ�-o{Kk3ɨQ��ROb
6��t�I1I����hA�#�4��l���HJ�K��@O�'�w�D��H�CUM�jF������[c�9�7�`r�1�G@�z֎y�
����-��_��5�ʼ�̾�|Hu�8���a��5��zt�h�A.������c�>�^XB�*?n�|�����kV���\X�f����tX3�����t����V�H�we.�����yy
����������L��C���G�؅+�"�̺��h��O�h8GT&l�h����jǔ,�3��ʁ���,�W�"����
V�/�:O��?\.<��=@ �Fx}qX�>��V$�*?v�*��>�)eO�S	�H�h��OY�&:� ;U���]ZT����W��� ��	�I[�����*{� 9�@������(G�ؚ��;�����$?��UO���\��0u4��$����~(j�Ӱl~'|��{ö������SF��+w��';�[���Ě�]䈥.f��f"��`�	T@�,	��K���879��Ge�\���*���w��A+󕜊P�&MG�]b�?����Fh�%/��%��"/=��Ntp�4էI�,��@�4�������������@��+F�?ZF�m��1�v���<o�t����\������g�(k��i�?G�z0�ba���1�(�Si�NB,��m����Nw������5?�#�_�pX�؅hi�u�����GI	��V3���d��S,z���K84jxp��\��$�!@��o�-�B}Syn��.y� �x!��bE��-��)&�A��$q��F���xf L� 'O+��`%�
����&,qGh�̨�*A}I�^�ٱ�w�����#Ů�=[B ��J�%���$PtO(LY�7L�����o��,���H~��t�N�����(+%���s��j$Yr��a���kj��#;�'�h ��~��r�5�ś��x���\N���Rk'Zi�@���5�c���y��;�q�M�]bWTB7����:靻3ݲ0,�b��m�P�n������/Gd�^�`-2E���Q0Kk�J��U%���&���WL�O�p ��SC�e1��BTcf�⬑u:@�L�B�s`\^39��<ʣ��	����+�u��-�C"��H��~`xL��G(	���b������YUX�4�:��t%��D�'��i�uc�1�&��d�w���Θ=�-:{��6�o`�t�*\V>�.5T�d�� ���4�'����N,k����Q� �F��-��o��������7jj[A�ϵ��[Ka��Ap/$Q���x�䧴�����q�tz��Ѓ�.�Jy_?{̀�}�b�<�<���z�F9{'�ŵ�b �L]hC6�`@�Ա�\�=��K����.�f��@r�seE]���� @ ��V��0ƃ�񫰩�U�$�)���N#@~f�1���c'�{��L�O�
Yn�gX$D���l�2
я��w([�\�<�ļ���Q�@�F
�$h9�rљ�~gCё���qҁ	.�|��O���.J����� "j_w�e���S@蘋I��'u����.%2٠�ݛ�9��K��2��b�L,B�hTݶ�fB�U�3j���TCd3�S��'�����i�����m�&3䇧�'��Z�&)t����H��=+s�1K�寴�0	� ��pِ�� �}x`�ekߝ�)��������~%�z���+s{�=ߏB��j{��5� ��>���c_�2�ˏ]*�]O�N
���T�@F�����չ!?.)}K�>J�������XU�B�W�y&�Z/$k���*C��u��WU�h���E������^���� ����O�,NQ_���9p�gpԣ��ẅK�T%�EȅrArxn���@a�8�X�5nd�5���SWj���!�7�,�P56��3��(�3<h�`"�6M?�vRd�f���ؔ�ƴԶ���z^AX��}��~����m+v��Y>|��@H���%C�J�Τ:�p�2�49���۽v�{�����\UȎ���d�C{�/�-���1#OS�������`�e�$`ɫP���H��#	�*?���e�����E����jm���r��5� h����	�.jS|�`�^��]{K���f���'W�DF�Ӯ;��_�	T"���I��p�@���c9;��iFoNҒa0o(�:_����o����s��-�����\�)j���X ��L��<�qɺ������Q�s^8�kϬ.혀/(De�^�0���wx��v�A2I۟�\B1w�0ԋ�D%G����8
8�w���oP�f�	o:�����DF��E\���㣟�˦M�:~��ۈ���⏴b�ܛ�a�7�x���+���5�I	�A_�7������Ӂ����Z��=����6�]�O2�E$��
<M�^V��V�������0�3�q�����<�卽x�u��ɼ$��&T�te�h;�B�8;����Q�*T�����l���5���N���U>i��2Sw��!�2��C_@ٺ�+��J�A�}�>�t"�K��L(�t�Ř͖�0����Cd�5>۱�i��!��g��t�����B!Pm��-���#ƀ(�PVqY�	.��.����L��4�.�p�12١"��c&��)�&([;�0�$����m�T��6re��$�y��Q ��@�c�{'���i���/�l���r�Ĕ�Z�@�%�E��(+�O<��S��E�_L@g�9�z/B����(�[�=�A�W�/c:4�*�	ߍC����j�Z�U���WM'�n�$é�'~�I�eAnIk���j̶�D���] �y��#�ͮ�-ڒ��W���E��,�3��#?IF��_��1�s]���[CB ��@S^���Y9��>+��������<��|�1#��	��?�7�X��[�gD�-Cbo������'mv�I���"	�K ϖ��9א����q 돸��i$C~xTߚ-D���p�.]�ʟW�w�p���h���A�UP��ɺ!��OL�<僴�V�����)�����>qL���QZ�3�R.�+��LZ�<�� �� �mYB����Š�,`�u���P$�����`?�����ع�%��
7ޯ�m���e�լD@�փj0L��A��a�ww�Y
��Y���`	��͉��8�Y�{5%�D�EJ�'��h�ή�P���ױ_=�t��J��8r�2a�D�8�ă#CYT��R{��&/ml$#�\�n����\z�Ԃ���O��Ҟ;Ց�LĲ`���e�t��Y�����'YH��N%a@��0�۠��m�F�{dab��)���B�	T�i\w-$ߘ�̗dͭ���}.����]�|��!�oX�
��ң[VϨ}��6�0|�1�$E�8�9��0�:�>�%%F�]����ĩ���\L}Bx��v-/x~��<l�R6an�_�'��@������̥\ܐ�_j���f�F�;��h�! ��xF�F S����L���197��7�cB������-�󥷖�ԢRV��]��-�k<ߓ��;~×wM��a�-_��<�ɶ8�ǵ�� ,w�p8�x�ɝV05a[���үQ��.�&�o���>����/I���ߝ_f�^O ^�w62��Ƙn�.�'c����j��w1�������89��
��8�do<R]�a#��� O�u䩸��3V������QK�0����ä�L7"��j��X��lz0{��u�Q�jD,\�̧����y��g ����M ���#���.��Ϲ{�3A��akJ;�e��	�}�(2�>j�9���mA��VCzƞ�����J�Q����dA�e��8k]e��ձGw�	�/>S�~Y�z��\T��pZ���v�BY�y<�fxg��X	�?{�[ɟ�v��2�"��ׂM14t��R��0d��Hr���^#��ę���%蜜�P	{m�g�K�< �m���7�����FL��aÉ]���؀�A`J�8좣z��Bntڹ��Sv�\g5�]�"�4�xv�Tܸ�!(�ͪukGO���+��Q:�9�Y?��sZ%$_��8�v��ےk��|4���6��~ֵǐBPR̯����Q���	���	*�#���7�� )J��/2�i
!�~(m�H��5�X�Գg�`B���$�o9���m�y�H�tb/;
�f��`ĻelG[�Y��X<+Z��ֱ���l���rk�l��#	�ԟK��If�T?Mx��j�Ǳ��D�3���(~��fW��{Z����#
Z=�־k�Y2�/3H,S����43B����@�O�#Gj�
h:n��*wq0G������{��<���lh�FB���O;�Q�z�C�#w;T������Zk�%R��9�Ǥ	*k�����>��L�Y��g�j���KOwL��~+#�����`�0�RGkV�処��?:����l��|,V�R�*N�~�d,�3�c�R#:�q$[>�7��x\��d���`jv%KVo\���Ax�J~\T臤�C�3�y��ۈ�v�/6�!Xχ��6� p��jj�T�I`��������Tn�����Y��Ѱ���C"'(����(G��g����N5p�-A�:Ӵ"�]��Ҍ�28�J�u]$�,c��6[[QO\۔�eқ�B{Ҙ6s����3\@ ��8���aS��)�;%V�VN�{scA�{g�D���D�ys�	R������K�U��X̓������S�̾
Y���Rا?r�Ѫ�Q�
YH�+0����i*:b�c�]�&�>�����:�"G,�V]}�s��X����?q7n�@���h��-��c��h�POw�2�9,�N�),�߷g�iC�4P.[9 �j���.��G1Gӎ�`Y����Y{G�na�P's��\��hb����Af��l$������`��JׇUv���w�g�}��C8B�׉N�[;g��gjI�0�c��%VV��G�Ҡ��0�ؽ��)�EȁUd�/���9�������k?��S!��uS�k�=H�����xJ͏���1�$�<�&�	��17�-�H��v:���&G�YQ�eP��ҿ|Sm������ &�c��l����&���)����6`6��w	q�` U������	.�
saX�� ��H=\�/s�x�S��K��2g9�k�Fq8iVKX�c �҇��s�όs�v<���kэY�k!�]P��蚭F�l%l�WY��M�E��Ss{ot��|�m�IY݀�g���,�~
ϗD���M-�3��|�uf��o���0�|�n�L���j����֮p��v�����9-&�g�o�f[�����a� ����Bvx��*`��GKf��l�)�7��	h��C%������o>a�y0c����-,�TRf[����-���v�ۦ�1?�QKaz���E�.��2$�o<a��?�xVw�4 8�	rr�:�,�^!�ltҳd��G��A��ǽ����#�	B ��y��a����9o\ڱ���+���b>o^f�a�%�t^xlԉ�Ü��x'B CTN�}��C
�Ƌ!��u�4���;��bV� ���2��u�+a]p!,1}9�I/s����ϱ��>��QW��%,��{0`�f�h�U�;,����UeҲ�{M	uE �S+�i=��f�]���{��Ѵ�MP����(�]P8+*8�$�"ȋt�R~�̔^�ך%���'9=_��䗊9�c�׷�'�z�6������.#�e���)��]�	A�ې v�L������[�ww�m�[�T&|IM+s �saN��S�D�-�.+��� y����ռC��s��ta; ��N��&�������H�B��E�v�Y#㸠��آa
��v	� ���Qq���pQ��f�qw;�S��Kn��lW<���;�WD���G(�D�eb�x6������ӛ���;��;	̦�H�6�Nc:����k�|`j��V�f��.��à��S�!p��t�Q�'ĶN�7?����N�'����>�WN����,:��m��j��Kr,��'!o�z�D�#��~Sƨ|w�et.����Y�AV�8��'���]�B���2�%Ct�l�?"�Ԯ�੟�D��[����Jx��ﭮO�	���7�I��n�ӱ�u��t�ȟ�d>T01��W&5 �K��'I��gA�t*ܱ6΅^�$�.�]��ݺ��-Y�C����!I��v��ǡ����&���}�ȕ�<���L�;��{T�O��N�i��?E���-˿����i�
�V�x^<�;#���.hԅw1ؠ'��#=9���3P���'����1��hD>��� �F.YUڹ"MN��k���(�a�'盕�D�_Փ�P|N�}:2s+
��IT�`w�����o��~L0�=�0f�hMH4&�u���0��>iE�S>e�,JT���h�s����j�J���dM�I|���G�р~��-|j�ʙ��S�I7�]�#�8�� ��~3�(����"O�3(��\�{c%���o��
nQ $����E`\<Re�|`4���lrg��Vz��ו̄[�ڌ.��B��S_���u	�s�>D�,4���ql�}�����Y⳨ʗV�����5��.�1K��9Q�'�Ѽad�f��5�Lq���t��S�l�W �BR�����|�y��Q<�*�IJ6H"�x��Ø4wԥ;1ĔZWqkt���w�~�}0j���6�kO��[�d�\Lg��7�(��ͤ�*�h��6�X��sЦ������5�/h/C���A=��eE{l�!Pp����"Y��V��W�
��K��ٔ��Hͳi��Ct�?��gZ�F]/swՋ^14��}2�$NpW&`@�uz>^;���4{�g��X�y�8�1�ݐ`D��� H�y��3A���Ʋ�)u㶭���r
�g���
p6J(�!dy_N�4ƺD���^:hU ^���V�~(�6�'g� �����7�6����صna��|�%�ދc�瘟B[�*���Q�^][�J����JOl�U���p��M6z��;���'�\'%�=(�I�c��q<��o�N�K�2��ז���"�0-]��N�"�x�kQn����'RW���i`	�I��f�1e�f�d6;d�Q_1��@Zb�n���W�e��Z4�#�fV�
���L�#;n���	r+�Yr�j�b=C��[�4Z�F`�{6G�h��Qq��l��I�o����	������_Gj(��C��ax�$�3I����~�D�':$���wv���r�Aǧ�I�"`bO����c]\?�U���].g�(�)6���\�y������x�EWn����nx9�[�!6b��~�
�g�o���*M;aT3���N�p��5�Z��7�J�G&���=b)��&�F5�ݦ�k���Xg���2��A"�\W�ԯ�P2dڦ���n����O����=则�Q�X��.^���ݩ�9@�͠E�;|���-a�,������"f���<�8!zk�-�,�q��k�.�Lù"��!�+�9}�y�Le	+<�#$�i`m��J�	A���!�Ue��:&���a�#�\!�S�l�%n���C
�3��*Z{U)[;d.�=����Hp2�����G&��ߔ�\������Tj+[�\���Nk���P�{J[����O�,K��l��G����C�D24��#V׋�؇˸�e#崉�ɋZ�����ּ��Q�ˤ@�H=���I���~P��w�d+y�.�v�R768�4����;�ZS4�tz��/#��~'���ی�������3B�/7L�;3��`w�wk���(z;�<뻈���|tH���
�yS\��4�E�72ތ�'�Ex��E����#yP?t�
kE:�T�����������o���Ζ���#�I��fU���,��6����Iեo �*���蘀�G�I9���WjOK)X����'��x��:�4Zc�8���.#.��j�o��PGb)<��֣�[�If�m�`��<m�8�/X3L� ()s�G��~�g�v�UZ�e��Pه	�%�h�4�����O��z�G!�FJ�;�-��@0�uF��A�Cwc"��9�ܴ��y�]<Uy��v�ar�G@n����y1�pީ�����]|g�,I�W�C^��E��\aX��>����vn؁�e ]MmLV6tYh�*	SE�bt��%H��Y���T��?��<x��'p���U#g���[KՂQB,āX��I��Bm��/7Y7�G�whw`�O������g����lN�8�b�l����+�=~��ԩ�b���O�
N0~F�ȗo!������.��U�Hi�gt�%-�{T͗��r*��'�E�WJ5���D3�/��/|UVQ9h���J�xVs��{�%� ��e/?!����K�v" F}o^^�]5MS-�Xah��l~�+�h��D��+c���7tͧ�p�p�dM�=�z�M!z��A�b�;��B��'W�ȁ)Ju�/;>��$���m�Ub;�����e�k�Z4Q��3a��g<�ϖo���L> �1pb^��d�f�$���c0[�/�	/�<>����)�r��p;{�~�߱��q��*�SF��4�����d�$G�yo�L�<�2,�?�)�6UT	B�G����j��u��|��K��yqW��T�j)���b/�	fp��R���zpP��xqo���D�)����}��ym�D�}�	��$��y��]�ж&�P9�M,�j��f����	���)П3]@�!�gD��^S*%��F�U'�4+�CC�-U{�V6y1���f!�Fm@Z�$w�ׂHN��g����П(Q�-kG�G� /����x���{�:��er���Agv4�)���_� n"���Y �-�D!Z>4�XRQ:������'LV��4�Y�؊FT�F���*^��}�8�[Q"���m{OҔB��۩�Ƹ�3fXIt�$p�W$rIY~@�ɀ+l����(Ⱦ����@��g��0(TWo��_���%�+2�Ÿi��T����q�׌�N%��̆�k�!��b3Bg�1t
#��_�mg�}j�U��/��Mi��q֠>���:7���E8������bO����ut��Cw.
��--�͵p[�	a��u!.��A�TOP��Ub������2)[���s�~ٱ6/��T=�T0�exl��#`�X�
�&�\�#
���	q���J�<��mnp<P꺴k<���=e��|$�cΈ��j�^e��1ߢ/��e&�<b�ഷ��r >����L7+v,�bx���
}����fܞì��jL֠7�>mO�K�N��pΑ-�IW�4��Y���g�2��A�����=�Շ��}���v�;�5��f�盯�;U��Ẁ���7��3H;�1ޤa!�p�to���=�

1�o���=?K��j��R������ʰ��Ӡ���~�4���#�����h���T��bM(�SF㘁���]>C�K�E�JmOXm�ah��1j2�ͻ��c�°����>�?�ik�x���M����r�W�b�<7}�}N7�\_�Y�h3"{[�x��f��O���y�o��.��g-؏�D�U���P�Kg�y)��7NO ��`Z�� ����tA��iL�z!�'vb9
TY%���H�:7U%XH�Է!01W��t a4�#���A�Y��4��;vX;K\��S�Lʢ�aƜ�60J�����a��lf���d%�Ę�*�S;��֒��끗H�N��?E�d��Aw�����>�hϳ&��"�, �Д��$����^���M�z��o�Շ�J���d�}c��X�}q���E泯ps�E:���pB�����3�н��^�f�������cw��Y`%z���a�$q�bՌ6�r7}l���	CVi{������c����6w�Q$�6ޑ���!a�֤!áW�Sr�NI?��#Fv#�Mgk�����A{�£M
�Vv�lEށ�,�+�ڸ���~[�r�T�9ޖ���CA��'3p:��J���R�G���.B�	����# ���~P���<Of��\�il`5�4�i�B�)�����Rij�9 r�c��)#FLp�8C�V7����ݣ��:��Q��"����O��t\�,Z~����Lyw�I�g�޻�u,��MG2{�j��%{	U�+��͉�$� 8:���`�Gº`�H��LR�P{΢�1��5�/4�#����9����М0!2�}ҘB6
ޯp,�t�F�q79;��y
K��cY����;�����U�g9a`m���n60we\F�9t����3�!I�a2G�g���7���m�J��D<rd�Si>�� �0��Q��F]��#"Y��V��P�� 1?B�@+��v��`[�����ߗd����撣���Q���J�7�!lŏ+�z��40�xM,
lO
�6Nՠ��niy�0�
GE���>�~��5�#��I����!���В�\Y�~��Z�9��D����J5�e��ڹ���Ks=<�DZA�8MJ)d�����"c�G}4Mi�%�����p���|bq��~�Q�at"6 ��O����F�-qq�/#��+&:ݗ�A�C�GjOg�(�K�� ��A4v`h`U.��$�i~`zs���#{�?�ؚ2�'��+���O����,x��d8n���K1C���n�K?��k������}���������&2Oa��#m�M݌�;��Sn�|�'*��!�޿��31/�φ)>�B08y�d~cnP3h���Q����wZ�Η���<V%� ��Q�����Z��>��J��~�� 	�7d��	�	�n��(oX�L/��-�m����� ˢ�`��U�Rj��.B����8ڞ0�w��t=�tN��Bl<%ö2͔�v�]b�{T�Ї��#�㒿ٷ�0ڃ�-Q�N���V���l�~V8�ê*��a�:6E3Vɒ�\C���#��$���5�ad��旬`��,�Hu��2��aM�R�<������\l�p���u���b�#�r��Ww �h�z��F�$�	+�7�n�X�=k�Lc�L83��de��ti�fE��=�;:ы������I�8xc���V8�����џ���n��<�}&����'���S#]ՠe���AW
�����,��Ƌ��nf٢��r��c�ldc���� ���yJ��=�z(��˜"����t1|��+����$�Y��g��L�"a�'Jq��T�C-?��r����lv�K*K�؁]o��}�몈k�����a˝�#>L�Eވ�%01�Z���h�0$Z���iMw�`)��R�F���Doa����^�Cn�-��p��i3 /ERL&W�ϛӹY�D�o�u�z}����	1��5��j�R��[�~�]���`"<p�{��(o9)�4M����n�؀�aP|��ͫ�K�gp><�����H�x�|�&6�/��B4N)-8���`�:��	a`�o	m𡭑P�u���`�����n�U�ߔ��6(
{}��+pG/i��@{^�:|e��{�� )��f�->��R������g���0��*�K������fX֒ʂ�~�w��2��m�`t�A"�m���߁�)7&�w��� ��C컗����k	n�.��9S�l�(m��}J��(�/��Gx^E��i&T䎈D���@���^$ �MAZ}�{i�	肸,9��\#M&���t��%w��,0/8�NO�\���{�V���E ?�Rj��(��[\S�%�B����qO��&�.�y����ދ��ʮ]�ڵہ�sK��d\y#0J�U	o�в��d�������z1�E���muyc6��U�A�di�n��%�<R�E�4cK�qڱ�W���q����`������;���GWh��穤ؑ��o��ɾ��&�_x�"wm^������|��I���=��T,�B�
P��G#�iJ֚sS�ˊ(n��zg Ym���<k�����ǘ(�>�.�+&zC�2��� ��¢�1��|k^^or�3���z&p�$��{��������ZBH�Mb$��3�a�d>o��j9�B��d������D)
�u}�N��q�P�ھ���A���c��dLM��x����7=���w&j܌?�Tk	v�i��鋄�d&����'yr��"�V�WB�H)��L"�8��·5.��؂>ܰ`�����F0uӆ1o�O�G�����t���g}���,�M#��V��Ĝ׹��JÞ���$���m��P���^D����狎ȗ���%�H7X��͝���E��;z�]�c�� �nX���#S��jP���I4Yː�Lt�c��^���m@�+���d;W��<����P7����%�{�ҳ�ĵq�g��*�����$�@��s3~MԐM���B.����K!���M	��\�� �H�k�r��yx�%�������4����+�A!ʳ�*���T��[��yޢo��D�W`I�ɇE\%)Ճ!����5G��Q�T:O�v����j<��B\��[�S����k��S4j�z%�(����lm��Rg삌0g��E4T8��i��¨Ca�m�.=�4nem.ΒF�������j�+Kr�����_�"j@�㨾l��
ˋ�f�*�$au�I����"�+�e,�&ݘ���U�u�� 6t��-}�Yŕh"
6�R����V��ž�2�	��"�/�]�f��{���[�q�MLk�)�Ho�5k��;$�в I�4r�-Jf��
��]���k�GL٭*5��\%�!�����	}��������� c��"j��8�j��0DO���ի*ƣ/��c�֐�XI5Y+T`�I|�6/ : o���3ݑ(B�C�@��b����U��/�n�W'�L�F�Қg�PH��V�}[/�$��Ζ��b�Ã@H�e�d(���TB:�!"wRu�ٵ1�h��GO�8�tqh 'd�Y��I<I��u>�p�u�QX.{�%����I�:A���UM�=$������*ڝC!u7t������������m��-�����n�F��q�K<v���b�����v�MS��p���Y���(rZx����jQ^>^M���VT��qW����!e����m�
�м�������H����Q��������9��R�/Ȳ�WG6�N��ĠQ�p~�\Rҷ�"f��\�\詴�z��N8V�S��#�14Zo���c�j�n�qP���߳�� �ޜTݙ�Y�ɥ�֒�����g7� �%D�C�.��`�ӎ���|�L�/K��������8Gŉ'dw]�Ŷ}.�Pg�!K�F�^Ѹ��U�{2ڗ��{�\*#�\����48H���ь�n-�*ş��W6���P��9�cř�^�M���9�t�rwP���C`jH���[�gH����g�y�b��k}*��	YY�Q��gBb7q��D|��I`�@��f���q��
��@~Wr#i��� \;3���(AS�{Jr�iD��X���Z�"g�l�2�?�+$�r{�߻V�N*����EN�]��[-�x�ɖ*)!F�{g���`^��:d��I�`(�H~bdg���t6j1Rt#m3Ld�8i*b3-Nw��6B7fo�ch
Bh�e8+w�L|�~���GR(X�{в�@�ww-��7��;6�?~`/ۂF1Uݯ���,_��[1�x�ÍE���[���y��ޖ�M��-���oS���o+~���G�w2��6�J�%"��ԍ�����b�CxN����ᘂC��r�W�=Iׄ�n��\�n�U�6�`�8L:���צ�UܩsKu^��`#�da[�x
_�7��'!��~ �]�5����~�Ⅲ�[в%k�a[[����,7hG�D\C�-�F���~d.{)���=���ﺕ쬯>A�&o��������3aϋ�ZM�dE�A�r�]��S�5����l���o�@=�=��J.�.�9��A��a���������*�I��DF��L����n����>�����:�*A�]��<�i�4T�:OK��\����Ia��]rbb`�,Ze�R�#��2��c1J/�'��!������7�ٻ�Cjo�_h��f4�����
逴X������>h��AkM/ �3)��ش�+e��5�n.w!�T3�`S���J�^�'�>�%����
��$g�Qn����[�*u���ؙ�!�:�YE
9���� LkA���jމˑ�d��<��B�m$���oڣ�5t"���7�H�nѷ,��ș-	OCi���`�G���%����F*�ۛ�mw������"a
s��[��r�v�o7B����p�8�N��Wʫ�R�j^���k�+����]G}���;����xV�\݅ي+��e�q*K?�ei��g`O$�5|C���ο��
����g�<P���y2��o��2��8x���Xۇ�ᆶf�y���\l��Z:�[-_^��#c����?�lmw�R��Ьp��ɏ�]�=[�$�gl��.'E����Q��	5`�KL� ���ن�Ｎ`0�I�5@r�ѹ)��U(�M��ƒ���QT�NNpB��9(�H�U���@��~
M��NK�\�p�Zc:4'���L�j�j2
�Z]�`0дiڄ1�d���#��IqS�Wh�g���5!��g���0��h�Y��	�N.J�)�DEx��G18(k�AGTrau6�al�GNJ���
q��dG���u�}�K^.�8�W�m�j���C����F/Z�A�L�RD'�Ϣ�Fy��R�e�D~cU��/8�r</�i@��98Nh����B��dqh���;�(�[<��K�j�� ]�I@�Q[?����0�Y��&c��j"Ԓ'�w3&D�
p��4�H2��K�MG!��g���7�ɰ\"C�A�Oԭ��kW2�_\���M�׵!�쾌M���;T�p�B�ڵ�fl�B�I�<�<de�x5[+�N��Ǻ�L'd��e���Qx�F8��ʗ��>���i�hqdU�}@Q�rd;�,b�,\��&OB#na���PˣPZ��)ҏ����_���4ߋ�����u���;�{#��w�g%כ�D�k�^G���8.�~XN��)A���Ȇz-���]Ee��+�����85���v��}��vJ�C�<���r.��"�JV�"���,���㴈(
~6��^�!U���	�u���iGQ7}��ߜ�قTNʦ��{��h�bU��O��� ��f:���
_�x�B�s�9"/��$�hڒ�엤��<g��jQ1!��'�\.�6QNhX����*���VJ&�Fy������GĲ`g�]Ǔ,�+���$bE�JVL��=dz�v�DoNQz) ,����H�4Ĉh��F����#�:M?�m�������K����r��'�|��,������� �C���{�˖�Ft�����'?��-��O
d���5�d���w���&�X��v�y���'�5l�ꔹ��T�T
���.�D��9SQ� @�O"�4^��ǽ
�}:� �V�"�5Vp�E���<X����͚�`% ��DI��	;�����
�16t�N�����y��/@�����*�~+%@̳��št�o�S��������>���\�nJ5���4f�̑�y�t`�W�9 GNܚ��i�b��^^�_^�t���m��d�
���l�_��f��h��X�z�Z�k��g���!j��zB����6�U�=z�HR�\�����9 )�����x��3̰��2�@9���w��"��Wɜ��3S��9�]0EW.E}�g�imY�gj�1\�hJ�D4��=
�!�����:�5?p��n�S��z��΂�O=内��2�����V<M���[@Q�jD�Pxb{���'{e���Ua��Tkr��z7�)nvHka�K�ȓ�漴~"B�>nA	cR��J�'6��)�|[�"��_�j�`���C�M��gW�R̥8�M!e�#��^��5+47rae�d�bd�9!1�,�����8a��R߅kD��7u�֡�j��9E�q	<�%b2�����
���J��0� �/)��}�� ,�߃6tP�U��<\9Dݩ��1���
�aǉ�����3!��N2m����(ґ��̇��oR���?�%H�*`�g�;/+����фÔ���K����u ���$��0�6�p( �����Z2q����=����^�O��9t:�1%�{�v���:��*bRr׃�ɺ�H~9�^�l�L����"I���i��ѫ���Aޘ3�T-�]�P��n����e���N;����ۿbhHl潍�3������t;'.��(��q�����{F�`�Q�����v���e��҇N8D�S�pu�|�K�	��d�^AOѵ�������N�봭�tI� �)+p���Z�g���a0/'���O&hGc��TZ�.��R�lLrG�=��A2
��k8E�^�b�X�y]qKO]�A�9TsXyģF�#�5UBn5<!���O�%U˳����74
�= 
:;���b�����{����\M�9O	�ރF�j8"�BH��c�־/�m|���у�i��qh[:�e�dm�����Dv�4������~���61���d�;�v��7�\���X�O�Ձ�2�f�:�z<b/����P�|���5@���7�2���x|x��A��!������؈�QH�hp�|n��K�,�9�-7�P?����� �XS�۵)�EPs@�6N9��T���{*	�5/Us-W��Ќ�t3�|[�:�ף>H��[K��`Y!��_��ȵ��Ct�J"!_@J[�'�]E��#���uT�G��w	������m��\Ra�V?��;�_��'+��ni���ө�)�>��3���7���+P��Z��lf�^W?m����hs��#������K2h1��#o]D�ᨍ�R�.C`�i�.Y��ʈ��^�����[(�+����w�L�\���Ŧ��xw��ͫ��u�c6�E��O
wX�[J"J�x(*D�	^��ٙGdC��D���&QO��#7�^J �!�V�GU�Ø�p�bNa١R/���1nCU[���
F�K��0ɇ��n�B,���#������$d�u�~�ݎ^cl�\+�W���:��GxcT�]�v["G��F���/q6��N���i�O�����Z�ބ��A��/�p�A�ˋ���v�:�U�q�Y\"�q�[�QK��a�ƶj���;��p����U�9��B��I�"�����/����*���\�>z��߄�wtd��i�A���y{���U�w$�c��ع�*Ԝ�7C&	�8����
���8(���K��-w:vn�z}�>����@%�h@���-UǕ��R�	�����7O�o�~��\.BfE������Q�Ce�*��V#֨��n�9Д����'@�Fۺ5jJ8G�}�r@l�#|�O�R��X/tu����!�m2]��ybs'M)TB/��CK�6B��n�-��P�¢�2��I<mG�09�,wҲkڤ�����'����l�5ޒ��w(��W����d�f37�/�aQ_��}��Q�h���(C-ϲ��ċx����5���{]��X�AR'Y���:Q�H|�"�K_��P�T/;ys�3��e+�Te�؝�k΋�h|�ZE���(==��h������%�Dv% wN��")V��AH$)����>��J����vnM�1�B�9Y�~�a|F�a�e,��}���BNː�3�Eᫀ[�7��Ҳ���+I�JC�+����\�!�#%�P{�7��6�w;hn���@�4l�"؞e.E|>�ra�k>{����l��X#/����%kR��BwFJ_�OX���������ᴣ�;pP����wٚ��F^�(��zkݺl�� z��y���<$����F���^�n�:[X����;�U*+ͯ�����#?����
i���s�[�X��ԫǖ�9X���a<���9������Kn�ݥS(m������eG������'r�c�|����l����3�.��,Bv{��7h 8���U	�!	��k�]po��5�$�b?���Pf/X׹�'ا*�l�Jý�e��9_��S�^׎0!���QYQv`[�1"��<���Z:64�K;^@�����T��v{͟>_l�&A�s���q)�hH,� �w���c��@����/{b��إp�xAE���aB	ܭ8]�Q�w��F?N��x��v�d�>��������p<f[��@u��io��d��+��Z�:x�p����N�������]�IQϸ˳�]�m�<m��[��zA9{:�7cG^���o��D�C@	��k,{�uQv����N�2�o���3#�	�i�c.�B�J��[:��8�śP4�p��x�#�lP<3)��+,Y�jJ$�t�l#�$�rC�;��C:��6�E��,IKc��I���'I���O�1V�=f�\O����fh-d��wJ��Z�]��w�"�,����%x����Y8D��Фv�wO�}@�:�y3^(h6wh�6�Du"��XU�b,S����r�+)@A���$`s�.��䇧,�j����+3M�7F�����c�|��Ojn��a�i7��U�����*G��b�oB^��OB0F����Qn��|LL-, ;���|��{v���Lg��\�ԍs{�<��T5�RN�B����z{g����|_�G�2��>���B_��^�(c[8Б�@�#�D),�18o�Ţ+郌��?9��;ʁƵ�o�(�fzq-a���z"���R�ߐ �^?��ԗ��~٨b,N���.r�(�b���S���U��� գ9�1CX�L����T�������\��[W�������r.�c�j2ة86���BHKԂ��)Opi�#7�sM*��LP�H߳�C�v
��)��>�v�M�~�f��a%kpS��@AS�K�J�G|��Y��HPk9A���v$,h��-u@}��䑲�~Gdf7З��W������>�VC&��[R0yQ'R�$��%&�)���u���痄� �}�kd(-�~ٕ�UD;�T3Ʈ��h��_���hɄ�D<�q�Ϛ_�H�b#��ZO����,'mv?�M"g��<Q��C�r�
�ʡ-F
�,֒e���^���̀@�Zbۺ�1��3f}�*F�q�����:&9h��{��_��"o�V�$����O7�M���sw�ӡ.+�@TϦ=��a#$��R�,瞆��XL��6���b9���_,��~��Ʊq��м��,����c�ô��&t��u'���ଡ଼�:ja��h��
"�2�4��ߞ.t��	�fw	_���h���m>�j̺(����qų$+�"����̖tm���әp�Q�Y�$��Ò�|�U���c�,�1" *@�rr���7������ӼJY�@m�޴�]�ʩ�͖��G-yr2�J�b~:w��h�Ӹ��_Yi���7�!7��>X�i�~g��d���Ѓp��V������3�jL��p������9�:~�p�
Z��8@r0謥�*LjYn�<7n��E<��K��8a\�g�%�P�Y�u�~RZ�@񭹹�q�ں<�NU�R�Hx�ФX��X۸���u�EO�y�WF�A܆]���v/"���)�����{ ��Kyء����qp^������ŉ��K��A3��D�
�������۹?��L'Z�h���O ,����x����O@pE�'4�ȱ�]c�w�	�Ρs+��z��_����J`$#�1�����_��g!��5��	C#��̆;U0����JWUy�@���DT�}&y?/Z��v9-�([
�w�wc^n���$��� [}ؤ�G%M�3z���M��"k���G6�pb:�	s��#uPyҌ�ұy��e�[�!o�` Gz��#k��ODz�4�y\��z�?X|���o�U�����E���<{�����2��^F�_]�}��/_����ihP��D�r�h��|gߝ!�V�5�����tb�xC���s���A��]b"�$�J�b��?�M���K���Z��[�@�Q�$��wO�����@�?e�	8L�4^�Z��T���g�C�P��$�%��3��Β�	׳
힁��KSfbM]����6�\�;�L�

���Y>P�P�­��}�W:�z.~3PK@�8j�ȷf��Y}�����X�@x*q"�9�X��_��D�ն����ǎ����G��h��ܩg�ť�y��P�����2�=��/#Έe�OK�!q���w����� �͜�Jz���1x�C7�ė��H�=���[��kq �.W�l*K���* �oM�'��%����=i��,H�A@$��)-����%�H_:4c��L3=G�l��d�9�o��P��Y+�t&8?W����I �:�;v#G�C�zҜ�sH����:�f9��U�J�����Ȱ豇\rs��C���S鶕߱r�'o�0�%��lZm���A<%��_�	ˈp"n%�`��l�<d�Y���Y�;�Ä�ˈ� 5;�	6F.m:Q�F�&�dWM'����R�Ok��Q�t�M�Q������n���"�	�.��]���1{�Çg�64F�����;'�^/��B�,�qMLb$<��8�dϕH�n[;i���L����3Y��"������m��w7y��\��}��o�,E�L�2�h�
P���"%��D�>5L�֕�V���o����OJ��&�u��D#1<�n[���;�D��G%[�Fɕ޾�o(P�M���4p�.Z�zb�ǜ�B��.�|}:G��8���J���$��Mv�?�!�G�\���T���4��{Q�Y8Y�#$|��pw���z��3[����#}�qHƣ�@��^]~����jE�@����Z�6���R�niԬ��t���;�Sx��7CK���g�����X9����ܟ��9@Z0�-�x��&`��Ƅ�����刧K�=��r+S�_�T(��@�xmW�VX�k�C�g���#��g��(~���ꢛ�g���!�9�|�)%K�Tf��
M7�P=�>��':�h�Qda�`�R6�cjÚ��+�1*ǥ�#�T���kD�i�asXj�c!Aj,QD7���Œs_'�Pυ�j�����,��Ki%x��(��_�����/��ZbS��X��bZ1&ZM��bྟL$�H!�!U�UΘ8���)U�B��9���Ө'H	���5�1Q�ad3�80�t2`u�����F\�����>~4�5P\)�����"'\~��c�<���\��������\�С P�=`Ӟ��:����Xn5'�"� p�(��|A���&*M�d�v�3P9�&)֕���H�TQl�2���P��e���ͪ9�m�;Hk|�F$qO���A-�ǭ��g���B\��l �o��>�t�d/r�U�D��ut���	�'�����*g\��gU�|�+ٗ�MM��p�H�MB��ȳv�;K鬡��،.ʼ[ .�
�=���7$)�O[I?�3��x�Ӂ�zdmb��@ ���?�R��u��y�:O{�/�G9������^���?.vl�I͖���N�a�r�;��6�m�]/G2��a�r�U�,�ꓵ��"D�
���͉C�[K����@ZƉ���&}F�0�8'�֩�lb^Ii�up�&E�3N�Ŝ8&�'Ƣ*;.���+Q�p{i�w Ƚѡ/�s���.�n� /��pS9�{�[,���~n}�
jr殶�U��:���`k,��lTc�2(O��y����W3�}� nZթ�+�	#
�z�e=�D��d�J���%7�I�� SH�߽:�X�;W�n:��Wx���K�HЏ�+�%�M�b�;��k�[IT���5�bK7��Wh�`j�%�ݹ;zq6��Z�m�������ڂ)yq�d	ҍ����Ù�Cs/,TW���*yv�Y��Vs��C_�	���V2y��p��EX�%����,��Z=��!� �9�i����iC��k\v���{�BT��N�L�����l�W��Z߰ب�ˑs�w�Ȓ�g����'"����Q�7M��d���㘭��f�����)A M&ü�帐Ψ����Q��x�;�n�0�{7y�㷝�<藕�)�RW�(����������R +��Dũ��;�h!UcՆ?�<:3WbP��P�c_�$p�Yf��@<���a�����GTіut4q����*����ނ[���3���@��<�����$b�u�%Y�hJ���9e��os��Kq2/�ƂK����_�Y�|�A��)}�f�,�!N��xI�P9փF�+���ZR_�<�� �m����+ǉ]��|����{3�sH�� ���Hq�;�j�v~�E����z�_�řꩱ,��wif����x�ˎ��6��Ĵ7�����J���<|���I�?_�׉�>ޔ�Oz���K���������(�k�N��B�Qʟ�"g������3�Cx��� �&�ݺ�kS;,qh��X$ l:�->KH֋�L����%��:����,�Zf��!���uz.�ic�2$�~C���s����r��ɏ�#�eڷm^	/�����tG)W�Muel{ߤ�6	��;��ܱ�N�;�èDm�eD��w�Ʋ�OkO���[/�i'x�9�Q�`�l%羦f`����4Pe�/~���R%�#��I�\��*�wh��*G�u�̹_&���R��ق��'��Ę��]���<�0�W11�}|bIo��@Y��^o���ݑם��'U��2�p�k�ks�(u|b�}�ؖՒ�'T%i�8�ۅg`�}�Z����]<BnqMu�Y�ϓ�v2��;���iF�.H�ہ*�7�ݿ�"�A'��v�7����^~�k�z>�s�U�Om����
+���b�=$*9 �m'��^��]��~����	ڙE]�3��� �������"4�J�(4���� ���5�c$Jԩ�_i�Đ�E*C�O{"J8R�U�x���U؝V���kk*��z�^tϸ�&���)������a��uw�z��3��ϛ����p�@�O���
���i �L�N;bg�!��j?�c.[�F~��{�����Q��ڈ��aF�2	��Q���tk��|�?�P$����\]i��ʟ�|�H� �l�2���%�\uG�"�P����C��x�Rߵ����|�h%�T֗��!��$�lA��,u�筜�O珖.n	�I�)D:���͈���� ��z�Y4�X�򵌑#��L�\ܧ�r��8�?��B".��Vc���8&Gq�!"��5w������?�����I��Y�h��C	�u�@|^�Zae��J���)��B�K|R���x1?�j.��]���.n�;@��[o:[���CZz
�ܹ@��Hv&-|Pk�P#r��zVGz�� ��[F�^�}Ʀ;e�%�Y��%�0�YJy����(i��<�1��Pw�	)[���D�7g?�����&�ɛ"[�f�4��dKQ_��'�B��1k^�؝ k��Eܼ<��}�d"}.b������IG��
nH�0�ړ��BÐ_`��ʾ`HcO�Fv?�¿Ga�ngF�;�OJ�������ZX�\_	|�i���c��X����wo�QӪ��T�n%0՚����b�"v���ܷw��=���N�隒���լm]���\�8ڛ���[�J0�!�}��>�s��=����~k7,Z��D����	�����˧�� ���X��|9a�|�y�a����
�U�H��2</�M4N$!�{��7}��q����:)_�ܵM-Ϋ���u?_���5�7�	K�0N���s<�8�Txx��>� >� ��������U�\�d��ATsX��~���f�߁�f������O���.�^Rp�$l�딻q�P��#��4aH��i�6�D��Q�ѿm�!~�"�*`W<�M�Y?b�-2r1���E�D8���F�z ��RnP���	�j����w�4W���~g����!�s��:|% ���8U�}�C��q�@9V����#%��:!Oy���J�B �4�8?�m�A!Θ��on�nѳ3�i���B��
���#t�:��WsD2�w��B%$
�A�Q��Q�[؝:��b��}b/
�y���myώ`���e��?��ض�W2��ƨ����Y��M��׶�t&�A'o�g~-Һ�AxT�f��/+����eX��b56��=X!;�u��q�dz
N�2=2��[��&�^�b
-;��P�G<s�4H���>��8�Ϻ�Mm��P��� �V�Oq ���C��6WRA-Cm�����$�l�Q�S��כ/k�a���-.v�. ���s�o��W�t4�nm��������)���Z�[�t�> �����⧦�4W�KO	F�n�g��T0�5E~���T�w�k��t��T���O�%6)�Z�"a��]�7倸'���7bŭh���^�*Q��!����##�,��p��O����M$+�W؇�~\׻��YY�u�\L���/�N���������H� jQ�s)cuv%�D2A�@�-����v�����d(��7���or�3;2B �\p�Uiλ�2&��Wg:�h�%$`*�ȁYni��N�\�e�1&��XRG�t>7���ЎoQH����W�0]�P
�!�Ʃ(���گ1ϖ~{��
ɪa	�o�n��9���Z��h/n�f���lHTQ��=��$0�
�5K��nan��%�x���¡r�_?<�1�Q�tQ�'O�^n�}�U=s��(��q����B��/w�K	XB$0���/�[S"�7�YD1��@t�-kMU9ŝ���0�E�`�naC�nR0�)�a�OC]��\�>��	@�%m�<��:P�'���NW6��N҈�Lpg�yV?^�ˬ�NU�e��	��[*�j�[���uKu=�����]�Y{�8e"8������ҹ9a9&(ߜ)��:B��>�ͼu���&R�:WF�vЫ�V*�(�z#�6O�cSۮ�{K�ђF�� ʦ:5��75HD|��=���q�������q��ж׃���ռJ���\��:}��nd��
�B�@�5�߉�>.*M�8�!T��p�+w1,����F3�uc��留���^����n�9�GBS*�n/@L���gu��2D�4��b�o�����u?����m�G���jh�?�谿�O���a����|�LXV�%��z��h.?�����FY�2%��.Z.�%<�Jz=���|�~��8����K3?($N��FP<l���2�<��>0�����47�'*߳/��u�{ƅr�!���)�"��?�zb."�t�?��#��$�-�6:��+Ʀ��\ӆL�D�͞�V/Z�%��:�'�W9}����X/��f0>��w��b����M��8&�B/�(�%!�M3�} J/��t:2���u����!�.�jM��o v���*��ͼ��'Y���n/)����G�����cp,B��կ4�������~&!�����zI9��!��x��dJ���6�#<�wA�T��qPY������(<���2�F-m�-�~"��K�o�̩����9���PȆ?ǭ�.z����^, þ�3L~�)~H8��Oy[���gU���ނ��(
����[BYx����9gb7�K8k,6��\a4�ʉN��̊b�r�C�7�[G��3�JS�#�����Mm���w�I3�T�V�6����h��� �˓�1J�cȮ��m���w���%�|�z7�j��ujD��P��ժ�5��u�qN�l\�# 6h���d�e3|]Ի2XU@�N]ӭ�5�&㪎d��bL{gu�l1���=�؏�'�rw/Ͽ��V����|��P� ����^����>�W���4���U`�B K�[J��9�c������4E6=$��c����g
��֜�đ�S��	�
ɓ;j��?�{#څ8d�]��5A���.��&�K���!�_J���OC�P]����]@0����gmUCh���Q[��R�;��s��p��8�����x�˨�<�U�;1aN����;>�i��9v���Y��-f�$������|���s"A��>0u��\�;[����W�?��x�2��e�`K�@���QL�d(c��V0�d0�f�e�y�{���)�L)����&8Z$����E&T�n��-Z�*� ��:7sb�Pn�Gy�
�_����e3��ɀ���T�$�3�ئG�D,� ɬ�[[f��K�F�;̑�}�#Ր�_o�<�f�4t�ȕ�;�ԑ�ޮ1as5l�-�i���Y��x,���p�M�A�D^��*���7�� ���r�Us|r٭�TX��˷����!#]���(�s�N�^���Z�g��E#�+�*+�Z9�e&v�����e~#.i�̇[͠Y�S��ͱ�uU�I��# ��O�lٟ�W98��xW=0��i�S��st��	)x�����r�<O+��+�s$-{���_M,�3�l��(�j{�_�;�0E��t�f�咭
����c멿��׼Z���I�|��l��E��C�F%�0xx������	A��r�B��]�j��9@�L����Js��#�B�@�MD�E�#줆�e����������yZb�3�j2����u�e�72Hd�8�0:�w�'S�F�s�}�����E�j��o���+a����`�*��e�Fg�VEh���.����*c|��;�Я���)΅�+x��+_�lE�Vm���+��Q�ܭ��`���0��ߏ2iM�0*X��ǭ�S{�ҢN�lǫ� �6��;��ҭ�#

���xM���(臤tpT���z�"gʮ�������ޓ1X�t�no���&�����N���Cr��+�=\�?�ݻ�ڽ~���0�c��eT�y�݃@)���?���Pr�'-`!s�����*~M[��ǊI9�ד��N�:t���|C�y�oMWO4)Ο�P�_�#TQ)B�=Xǖ=�r�;[�z�K r�	��JI4�s��F*�Dr*��9E�Dmy���X�-b�r��|nٚg��� 4�4U	� aw�����69��jF�s�q��G!�&c�f��.Ẻ�㒠�攏e�ؙp�~�h�8��f���55�����Ҁ��&�Si#�	G�f�m@��G�dv���!0>�t?Qq�n�ό��3Ca���Ҩr/�;�=��{�q�򾢥x�-Ӧ��f����Q,�CBBi�%|���b ��CV�uZD�A� #c�.`\��!+�h�л|�����p˯�V�CF�I3��S�|[�	��g[�����Ehx �<P2�S	j�rgƃ=%.��a�Gԉep���'t����r����  \>!�_��Pw��H� ��{�mO���2|��SKMQ��+1@l�e��E&����2
��a���$����W?:I�s��@X@�;�5��
A�11�&�]e�ѳ�_#s�c���������!)9�z�EXZj㖄ߦ�?�(���R`�G�ê]N�9��ɽ�>�@���:�y;r�2�H����*Ai�E�L�0�+s���QGvd����yDN-?���u�N"L�N�5�.z�֛�OHwɋS�N)c�a��ӄ/z�=Ā:wx��#��	1��ċ'H ��.����|B3Gk+A:�$�^��K<�1�vI�T�E��X���ϗP=�4�T���8��hj8]�$wj&�ڻ�"\Ր��-xbZh>�&���H@�6��F��Β�P���՜�����>r�!l�`]���h` �U�Z�u�\bgO*�2p6H�Q6d���v��K{v��cJݟ��ѥ���zקթsKCB��4w>�	��-�����H2x�o�<���`v�v��cV�&=%b��K�l���)���[�iJ��] 
azV:bM/�Kv�̎�;�I����P�>؟������_��:%&@#	[�A_��^����MS���[�1��7��9��^���^�U��:�ˆ˻���Y�q/�~"���[��?Hm~��P<Kp�A�;rvQD�M���o@���+�¹��j��i[��ɋ��8�j���OM��f�9[|>=��V���:�w�|b���{���H������Cŀ�-}/9�tj��q>������?p��G�ji��~���$ö�ϰ������1�`	[�26�
3U3��%zV�y� 9���7� z�F $�l����,�!�*���л¢��V�����k����(���@Rx��AѦ�ND�k?�8��n|�z��|WlR❴���rV9���w	}�p�����yTbȦ��C���v ���uT�E�["�)��5Y~��0K�Z0p�;D����WH�l�7� m� �
�{:$��A�h;��>����n�e�D"�(��qsg�@�s~��0F\�,���{�ʪ,)�&v��ɲ_q7�)�p^����1���gS�7�sKI*�ԑg��m��Zc���b\z��^Kl��;`���3)��Fc�Uhe�k�C1v��I·[���!�oL�p����'��LǮ�����}���p���o�*�u�]�����꾨g�1�Az@W^����iT;o6 |��@�KR5Ql45�S���8�\�H9��7΃�m�m��X��:c���&�̲�%dlfq�⇄����T�-��N��iy1D-��&���/��J���	r�|��BO�j~TQ6+ 
�䅑Gr�,%,,+�Ul~d�HI�R���3�q_ Ѳ�k+��_�c�ln~�� �*��_;L�,6�k�قZ�G%�v`�qBh�`�ڀ瞧��ԩ�I@� O�1uk�^���ӯ�}g��bp� ����n2�W'�~��1���Y��U�p�TϸS��/�ʖi[0��2�H8�ߚ)�7o�\v�F�C�*7!w��d$t�hh%��Bz6D/3�g�-Cd(�~gJN(��WPR�1b�����g�۠p�y�)V�0e9X�)�n܋�cL��.E�I�$|�e�&����v2δ�j� o�hѶU�UHFC��q w ؔ*�������؟L(e�
zwr*�Wm��_����ױ��#�O�P��O���C��ܨ���'�����/j巁��=���kZ\6�/}b�b�Dܫ�Y���X�� %O�SJ�o)a]�:{��m	���E�ٝ��i��|��tT(V:qzg�X����h̷���qmy��Xͪb���������N����[���S��<���΍ql�n@5`Ǚo� =��+�YxT����$_�=q6��l�-�7ٞ��������1
��gp���_��>�j���C�����w�Y�j�>��M���Xf#�U^��x�8_!���u��r�I�3W�%ǁ�M�A��p ��{�'9���u�%��RIu_���OvU��j�T�E(v26�̔����No����:�1��Lz9MSQ�½:����ÆC#�]�yzӔ��xq��B��-�L��o��M�5k�SU:eˉ��s\��;2b��Gc\]~�U#٘D��d��e��7!P��͚.,N��	����	z�"G<�x���"��O5 �h���u�iu�+>JG�2q��f�������a�x�e�iw���������}��Eq_�5��/u[��E?]]�-D���vf&5a�u���_��:�І���­sQG��_��#m,\y!}�z}���z��3l�?���7'
h���� p��������	�o�e�=�H&2� Ep����zX�k�����3 �o�N<���|�L��%�7xW��Qv���@���U?t�IW�G�#����A��C�"I����-���w�DFJw�X���@@��%��3��G��B��43�*���,�|z��q���ƈ�E.��i�T���7����>}��Յ�]�<w��{�����2�y},�~Z�#�{�L����2���/;�8Z
�G�}%oOj�T����|Â5L�m����h@K@Ŕ�Kc��0�<���>�%��D�z��(�����[=",�5h�`[��"�wG�Σ��2_��X�Iу��mL�+N��`��G#���k��r��������,R�iey���r�s_ɚ��E�x���uq9�I!��Eci�Sqkx63:Ha=� ,��5���w��Uͪ$�M$��,�3q[6ryOZh���"�cfd\��^{$={;�3S���M�?ۍƵ�۔t�/�I�z�X�j���(�eZ�'�Be+�l�H�v�niJ  /����R��>�;�r�g��Z.ݮ��ld�z����چ�'s�OM-*��R`d.���uΤ�P��0�e��f4c���1{>c��ܩ�����d��FQ6{�Q������MS3�(�M�����	���z�5/T�p�v�&6W	l�w�ĔSk��P�AxZE��
.�x;�sjZ��C��o�����4�y�OǢ�^n���F�"@`�iz�u�zx��V�����0��n&v�/�z�&�t��R�[�I���x0Ub����H���d�N��v����&��1{$gal�X��@vv�"J�l�LHkٲV!8�VQ=�,�ä��	}1� ��q.ɹ���("�i������Gq]�:Y���gJ+��1BS�0i�=zʤՅ'���޷U5�>���y��ׁ�'u5XB�ʅ��Q�n`��^ꜙO�ь���9�E3&���$w��'o���|X�WA��Q{*	�PO�[�.8L7g"�ln�)�]I� ���*�C ���A���a�
N#����������&/Y��%e�0ic濐S=��ؠD�:H���o�c���-����RB��#�X�X�ܜ�Z��l*������Ｗ�X͸�� �?"�y���7�yx�� �m�ʑ�V����(���Z�����חɇ��y?��]��"�B�$qT۶���I=v�d���F�NI���~��Y)�DpĞ�W}��S�Xv�:(�|��K�ZZ��:[Ъ�|.e�O�I`ro`+��B �,%���V�r9nd�� i�IE��[*��,�J���A7r�I�h �i_�g
 ��/:�㟗E�����ЗY0&��!'ZWPT��_5߁~fk6$%��4���M'W�<G����ހԓ(6�[P615�Q����>�����
v�8p�d�}��4�2W�Oh�K��(������@ǜm��$��.)�y%�i�����a<����/��/g��&/4�O_5F5[S�#�@�L"I��n�R���@��<���XǛ������w�>��P�U応���0����>�M�U~�Ji���ݫ*�kt�
��i�Azy�94��0A|\#��-%�f�������a,F���~��a �{U_�2h�ӕ�+J<�M����R�1Q��Q�����?���4��8w��i�FG=@L���U���]�L����z��@���;a��R?�����s&��q(�Ss�� �m��p���'��Y��Đ�����kd��.<n����_��p�8@FKN⧋��%��v����d��3�ǜ������j2�G�f9����]J�,�|Z�S�,����h��|�>0�5��l���9�+�A�E��8�}B�������o�F����F+��_����V��ъL:��g���ݡ���^�ūT�����"�e\�s�]ٝ6��"�7��R��*���pRS�^w�t�
������C+�]r������K�����0���������7��>�C%V�+����c��G���A��H���-��w��SI��xh`�S�*����b�ñi���qg*�*�� 1ap#K�.����{Bu���2q��L������͊%�����"q-���]�ɚ��1뛻r���'��b���k�'�&�����V��5��}�<�=�o�	:c<���R;�򙠈y���7�����	E@���,�4�g�l`֋ۇ�k͐��w���ޝ6sd��w��7��Lb��
Q��)>�!�~�v�ev�u��̡;��Ī�>2u��P�uCE�$���r/O�vr$��l�Le`k��+!��)������;��60W��YT]��HL�B���(�����aT��̅��򘦚����:I����7v~M�zs꟤7]�Sb��)���vDS�@ d��PB��+��h�O�!�%N)�D��=��}��+�+��=bm6Q֖�W6Oio{�
1?�k�S�k�W�8	��U���R�yb�f��������͎DMd���'>3Q�o}DP=2`���K{v}fޱx�s�L���xtI�l�(�|��-+]tYK�J�Z�T����d!��ӕ�_��)ه��3�3�������=%J1�s+v���Uۗ�)���a<Ђ��Z1@����ܳ�x�~�i�<Ѓb2J��
�%ϣܛ���#�4����"w�Yt��k	���8)��YN��YP�c1�\P��+y��Ս���<ʥФ�����0�8j=�V����n��tJ��4�c�zߗa���C���mq�ŵZWad��Fcb�_${�)�|-$��s�PAꅟҮAk���ZT/S.�TZ��PA�h�º꺞}+*)P�Q��䩦���w?s�ٹR��;t͎�ƶ(7��^ƴ8�\Ef���Y���¾� �s�x�;��%�X�7Hp��x�r��U-(����~\m�u�#�d�-���l�o�g�O�4۱�����K(p~�f�T��Wn6K��	���g���0���<��o\8��>$ɼ�sA1�������,md�1F�vy���u@c؊�M�̔�3���P�Ϯ�V���l��6�ɉ��ۑp6W����dl§?+�[�:�IG���"fvR[`:�1����̞�<��y���׉5d=��nu�:�*t@��y�����~%.��R���|��^�8zy�N��Ո܈�Y�C5H�{?}ٝ���6F9� �x.γrs�����Hѡ�pH���&�[`����@�C��sd��
 ��J�
IO' ��H����Ot@_]6�]1�&
�n����<��/�!��'G���#'0W�֩��H���س�w�|ν�8c�#���1����N�L6gI�۔�u�����{#������f�TU�ɡ'QFY���Q>�eϤ�cE2i<�'�3���S��)��-�;@�DݩOf��r��Q欤v"�c���\Tc�bБ�VE:ti��$x�'�;���s�P?�h�R�����J�I�c_IO�!�a��R�<��,��H�RX�c� �(�2��B�g|����uѓ �,�vb���ڟ]�dl����>�^�N��x�D�+����Y���z�@�=����L�sjH3� �:%�GpG��*��4��r��=ST��:�Z�oP#&��6B�Ȗ2rr�UBN��B��_�ϕ��������
�aYI����#�w�Ak�"4�u��g��z_�BU�G�W�jys�U����Ø��1Y���Y��\ȱ�m'k��[�?r���!{hX{�����SbI�7�;�j�j���{�����J����X''b?�g� �l��2l��q������g�{l�l[�u_)����_�'��f/��U��s�v�|dKL�2��r�(dh�-�v!䏿H��X�����3�Y�X�XA�e�o�����4�#�pL�)A�;!�ls2]���������^U���[s�1?/B�
VB\��z+4��?�P0��*�"� ޏ5��*���V��I(ʡ�;u^J����nw- ��-B�c�����ev
���5۰�ß���AI��H���Ú�`#JC���~��~uA�-V�Ǜq4�/f	(XUYv�	1����Ql3"Ӣ���	����S���f*r���e��+f;V95=	<���Q���opD_[9�'. ,�����!�f�Eɛ�]K�!�HCIv-�T̐�Ê/��U%����*��:�&T��y�W/r�E��#�U���d�������kmN�ҏ������.BRX5('����rHU(U+����'��$����&�?�&4�H���t�#����l<�d�Q�Ï%>I�붒��-�u`ۍ�?�`ྲ��.%���u�t�Ʌ�*��	���T�X��WJ�y�*����,��e�����m���ⵣ�2�rP]K�#�~����~��̧x�N����hbTq8��XO���9ժO�M?�O���G�������D�������̀�+��H2@k��8��\_I'���E�&}���¡=_w[���3EƉU�9�!"��(U���H�d��P4Ĺ�Ip�����K�	+;���~^�r�tݯ�|�c�kl[O�^��h�r$ݠu�	R�b�x��znU�~WE'g$G�Zn�QT��O�a�5�F8aO�9�]�a%.l�֟���,��Tu֘�I�kM�[��߯����W�J�m� |75G+$�2��ME�범vJB�%�ʀ�iψ�D;��#�<��o��:�,�.~ɝ�&�?܄�����Т���B��n�n@��K��:Q��!���\p���H�|	���/�T���^��<��4��8����Z~�?�톴��<��d@G�̆Q5��L`��g8�|���Yc?�*�!�TR�۟�ܝ��b7OB��6"�*M����Q)zF��������Ґ��V:1"���Vfk �(1ײ��DOhot*&�;Q���V�O�viHJA&��-`P7/fv�6�IB�Z;�Β�w��V�;�����Bർw�ǁ�!J=�ۑ# �����,)�Nt�f�d����k�<4�`H��Beà;Tp�h���\�o��ťM.U^��!�u��T ���O��Pӱҙ���q�=�%R��޲MQ\���?�k��G� ��P�z<喉Ƞ�h����˫�u�v��Lc�7D.R4�	+�3��8y�5P���I��ˬ�Tm�G7�2������02>�����6�oD�l�"���m=q�H铡`�f�-.���c�۩�ƅ��KZ��]����n/���V��=��º�a�`� �v��nw�Я���M�ޙ��AF���8�ɚ����߬�6��O�w��cY<(T�L�o����G�6O�=AmW�XI���P-�s_[�Ч�n`�[�= P,�%������j�˛E
@h@�뜉C����Kv+��A�HĆ
��ɷ�'��FFm��v�"o`DxV}_y��$)�Z����=�m=�p�?C����Ȃy��_'�;�cN�I8���I��I�������a:���p�E�ɠs$��	��  �����9�t\E�xl}���Dd���鳌��h�k��9�����A�K]!W����)����d�-�I准
��7��t����pk�L�_0�o�����	x��XNVY��������[s�:��L �/~����`�,-�aN��~[�\�E���Q��U������iu���0���0[-F`[7<��a�z i��L)��%���cB�I7@M��[�˥W��$�ѽ�'�P��C��!��f\П�M�l�7_,�A߆�9�s�����ٖVI�m��>��U(��[�E_b�J��J���'6���>��{��2�{�ެ��W #���l��P_Ҡ��_MG��G��G,[r��C�n��4\JQ���/,a*�E��W�D�*������w$��M#��5�� �F�
�ѴA6]�g���G�-�M�͞��$%�S
�Hq�O{�"�ʥY�b8�H����j��q����NH��&1Mg�y2|�N��	y����|Z�(]�O"��2�t�\?1�fY��{�5���W��O�ʞh����${9 ��D�Cl��Ī��\?7�(r�LD���
[ͬ�Φ���~�N9/�)�^��{�ڭ�`��l���]�O~�s6!�'P��.����/>���:���sWa���1ڄ�7�KpRB���9��TÓ�5m7�_?�$��ΝYW�~�� 6P�II�5&#�:/,�֩�Ί�F�S���z����V��ԡ@aM;O����҄k�%�|�j�H����(�]f���%f��;�e���U&$n%�JD1_��Dػ�]G;x�<m-"n�\ƃ��W�����,�A��Y�#��v���W�/i6jHCy�AM���IJ!�^A���bj�>ݍ4��pxkW#9O"��0^� ���2��Q2���x�Z+�)E-;v<��)�s,��z�N���:��������ɟW�r78wR<s��9�Π��B���:�Gb��B�͢0 �,�p<�$���Q�	$A,WF�bΎ�>ƍ\�����;�O!)�w|�>�#�]5] �ې����  E௽bU� �?T�n|EP��F�Ȑ�<a$Q��8���%4���Z�!���<��'p�/�JU�'��y�ߥ�$�ԗ�̯�aCȓ���R�����RO�{Vɫ�+.à��Óqt���p��g�$¿tؕ�^cQW�J;�x|VI_�6�$a,k��� �ol�i�F2�*t�7
�]�����N��ջ���PDa�!O s�x#��ӯXYm�i��ŠO��%�F60(~Q��C���- {\ݨ��`�:m�)d�}0;XƩO{���Xu~A�4y[��~Ќ�q`&]���F9N�j'���!zF:ja~(>dT]nYRk�5P�mѪ� 3)�rG��u�|�dzxoc�<at�f�[�_g��.���>h1f��{����Pwz��H��-�bkBv�|k�rj�����nL6���D ��L+���Oo�̭STLt�A�/,D��ݢ�&�2'��V���g��C��5��S��jr|�����)Rѽh�w�K���=�ǁ��+[>;�%d�/��Z�i��6��m�JP~��G4�VI�~
n��Cz�~��Su���u���`��\��Zy�'@eJ�����F"��c�{i5t QQ�̓�W���UU6�>�w�U��,��w�t\��}� @�c瘌�|�8��}�[�GDD�i@g�*�T3Cb�:Uq�z�Ȼ5ȪfG�wc�2<�w2����G�J�jV�8�	�E4t*����]��mĚ8�A�)uAk��s�i_�/�hWy�<YX�^���4z��n�m�f�3fA)4�����f�'uwj4���/�SG����(͚ȼ�i��-g�5d�	�O��B������p�ĕ8��ܑ_�^�M���PC���$�3��MGّQ<�6�v4�A����ݸ[R��� ������57������E�b��J�Jd�&��O�0�4g�W�̀�'�1)�j��<hp����^HlŒ���:�UDȊ�B=5����=���#�x��P`w��5^���N-ɜ<���"�z���8α[����p�ģ[F�S	��3��˭��MT������7ޣ�i�p���9�	I�����XQE�g&_v�Ȥ썷��#~�gM��)@�
�%]�%Ҷ�LvM� sc~=�GN�Z����=M�ց?����嶲Ѥ G	�&�,�g!�|Pz�i�y�I���X{��(>'W�b��o��2�ΟC$˫6�+���D@2?�Đ:����qY9eVc��� G��'8��F�b.����t����{eݫ;�#g;sȅ}a���Ă�� c�ǔbO~[fA�@����1�@���h�7�Y��7ڲhۯ��`�T��	{�cc�����+�m���g��&D��waeJ�5���p�V��ؠ$߉[�vm�6���q��s�(���kY��T�)��I5�e��PW��j�?#���]�ş�����1~�YNy8?��%P��4�ǯ#v�<����	�.�_C�WψV�w��{�*�̪=��r���J���M�U̲�9Iם��969 O�۫ϭd����N�Q~[�D����Sl��h	���3tg�jf�b¥���le#]��AIp���^⻒"�
7M�/��!����T8�
�W̴6�lw=y{;�o뺉겎���C�X�+#I��B#9���Z\U�f�ö��8��6���Q��5Uf%\nrtT v�L ��&d�п乷�ғ�^p)t�c1:��c7�4�������@��n���%��;�ĺ�G�Ĺӛ�l]ErU|��[��E�MܤƊ�1or��&aZ��ˇ�Tì1߆ߋS{A+VauJwe�0V�Ͷ:�t�n�8�
��L�= ~�i�����cm5��ۛn��U)�{�����Y(:�CpY	��8���f!s�c�-K�ӛ�Q-�:c�xiC��ʦ.z+e(���z%,z��Q#*-�&u�pO���\O��=C	�Q$��gys�T�DԔ#?�k�@^vf��͙�x�h]�h Υ*��s�?�ܔ�i�Ӥ���	x>e�0'&�}W�
�r�T;X�W����:��I�DA�)��<��I~֚{L>\����Z~��W�6��"dH�K%@o��I��`�iG�+F���m��ߨ��zG��)�����mwS&\�l��(�Xx��$_����D��4d��f
�b�c*صhHDV�s��I�
�:i_��n~l.�%��&��;h��$���O�������}�q����qIT��2\Lm�\���"�)�UA˰�a����ͳ;hO����Py�M%�oV������a�e̸�'��5ڔ%�1I��׏	�۰��	�D;�ڨ�.� �m�=:���q8ZN$1��tX�ѢI'��mԣ7���lf�i�#@��f�M������+^meف�Ð.���G�ڜξ2��+����1�!RIҹ	~���H$�,�4N�æ'ฺ=��MA��x�4��hC��pp��Xi���r��7=EC�js:��<r�tԍ��(�y�����(hbh|+�߆*6i݂M�y�p���'��@"�xES��V��BO�� c�}����]�&����o���}$��J�w��t94��m�gIف�P����Am�d�_p�E��PW��e��N|�x�Q��yL���;|���R�$����i)��S�+�����`�3�f��ƛ�=�2A��O�yD�:�r��T��՜��N �j\��Ny��^�zI�D˕�$�%;�cF�xJ�f
�ɚ� ��N��Z���3�Y��K��0i�>�rDc� �Nδ��e�G]��P!��y��C�c�� a`��5@�cP4��D��,7<�{���J6W�� � $6�"�}a�	f4�D���,��i;*G=R�րK�Ʊ��0��h��q��j�LS�cu�M�����V!!|ȓ[����v	�J�(�-"��in��|�'��ŲsU6�Jzxv�H�o	]M$7>�:$��S����ܔ"*&smۈr�X�Wm���zK%�����������~��}6|���P&�9�(��}�;5=�ǋ���:0Ӗ+����Ԗġ�/��K��S�j4&(����zZ��Ex	�?��`a�>Ҷ{�z�e�#(���Z��"g$��d_E�aQ01}���P�����֨ZmX�hb9jVD�=���'�9�*�n??�1���$)�X���o��RY ��=���3�L+��N��m�9�t����;1��c���%���\�j�{�1e?��r��󾖖�$�TR�������[\=_�9dz���:���=rL��]�«����\��R�-�w��R� �D,�Z�|(���~%�J��H�Y�U��޴���R�8�̗mUL���̅�v��4ye2��h� Z<���o���(m	xjx�8��U�H��d�[rJ�>��K{��|������<=؁�-<���
}s���]~/8��?������:���c<6��n�t&��l�k�'7�{��1��?���Ih�Y��S��vҾZDO�u�������7�h��*���n!��s�d���{7]f��Yҙ�/��.F'J����/3�Ǥ�{���&�����^��^���V�Iq��if�f��r�eq�hdWO�e,��2x�ˍ��?H-�*��$�f�~C�5��H~���М1QNQ�OC�%�2o�~/_y4�
�x�2z��*�����an���qLp[ ҧ���+�]�6��*^�6��y���O;��_�D��\��|y$Tg^1m�!�Ik�{@��H��Z�����T���`�?%�
�\�RW���bsQ�MZ5:����"�`�㺦�q���\/��d>R��8���aWw~7�B�\�0�R\�Au��.%�tP.9f��+���ը��50岿�#�F�U�ޔ�U�?���Т��]`7�����b��5��ph�� Xt�^0 5,-���]zF�v:C�=�U^�+�[O;7?NYa?G1
*�ר+��ݟ��Y����R��v���S1=�%���e��3����h#���De�F(UX�@�	�+7'9����Z�'b��#"o�H�_�EC냓l�*9Q=XgB1݇g�L��@MƓ�~PtQ����<lأ�l���1Q�Ι%b,2�XN-���ј�#�9(���4 .�?k��Ƅ�7��h=~A?�yIq�oY}��e_�������R-=�#���b�H�u�����YxE�Z9�����\*ڰ��W��j�3��?�_�cQC�L{�٧���&Ȳ��^�Z��sH����V#����쭁Th�y�$&��5	φr�G$�y�I�b�H��;/��~��ǅ����V�_܀��D�)���&č���ͨj��h��fA�c����邭?��?�!W���WY�7��z|�g��c�@�"�Ȍ�����0�d��dqq�2]Is1�Ű^�֭՜����� ���W���)��i���h�k6e� �9{F�d�ET-���e��r�?��5A�S�O��}%�gW�f��})����\B��U�1��J^��jrlm���ȑ�Td��&�%Dz�,�\/�d pP�KV�a�����{�̕��50���O�{«I��e�6�=���C޾��߉�&Qzmk���������Or��=���>{���)���QE�Sx��֜	�W�9��uܢ�|ӧ���6�����kl(s����,R�*z<�A��]��W�m���`�ʐ�z߰N�>Y�GřӀ �BȴyBW� ؕ�͆�Ո���VN*�0������V�)s0xQ��zȣ��ܙ��g��_�{�)V�KS�ra��)�G�bmߔsa>xd�RN��G�T��Y��7p\�~���G��$�F&�����v�u?��@,d���3&�MJ#���oGb����^��|�_�P�E�)�n̉�y�����fg�XY�Sf���u��l�K�����R?���0��%�Z n��¯vN���Hg%\��R͠��r���z�4�O*��G�"���f�俞�?1��"E<��g�#���S���xZU���ez��~U��[0�	~J/����Ss�`��tA*fh4
�A���k۔u-Y���E۸&��Z��|�{���i�Oy�Oߚ��S*�?jW���r/m�ܞ\E.�90��-�Kn����fe2'���/�pYm�g�03�p�ڡ�gF�����x[��M��梯Sw
�(�؇���ړ��FtC��ϼ���se����|R���k�&߼tr�Y5�ZN7�����Q��+�pQ�Ҷ���Um;�M��u�e�����{x��%S*���C���@�ڋ!�1*�'�o|ۑ���k�~��X?ٶq��*��(v����~{1*�Mު���4<��H'& 	�~P��>љ6e<�N�2����&�u1�}�x���\,}Lb������Utg�D
��9'��F�!���J���KG��'�nX2�~��0�K]�¥�ߋ��)x��f��&�0�ZwX�l��<�����E~��6�h��+=�<Q�u��~��"�wԐSD��#5B͡�������p�g�|��ō�8��7H�|���]��a��39tᲜ����7���)�[/�]�1��s!�8]#��d�v�K�;���_��;C+�m=}�,�Q(:��0�hW8�"���./k�
]�v���o��k���%H��7ٚs·9T���:͗4�z����x���.�dz4���ޫ��[w�a���,���U��H@��L#	�*N�_��w���ȏ�|.�ȟ�����C(pVY��IS��`��vq亘�=�`��?՛���`a�=sӴ\ݸO�D`m�0{PS"�7�+�͌��ɤ��S�w�eA,m�4j������`p"p���LW�����:�4v保�	C'��s8�R]��	R%3=ʥ��Dƒ�4z���9�&�N3M&�]�����d�q��rsW�B�����S^ʤE���]�mk��[���!�6�`���LG2XkUD��`������DB��F�S�7hN��7�|��{��Q��x�6�k���m��:g��J�(@ڱ��g��+���M���-��n�˛�洀ճ.k�η�6l8�.�Vy��Yg�8x�����0�%�	25��^��h��1%�"z|���x��8N�cTP�G��P#KSilp�y����wg�]뜉$DJNh�W�ȝ(\0ؐč*��H�y
�L�������E�mr��>�<:��>�D�ԩ��@�H�y*
�:�]����$��І�p��ߊ�圆&��ŝ������,���S�=	�9���ߙ�N�\4�'�aU��+nZ�4s;������.�y�V��F?��&��lGr�\�9,�gcS�$\c�m�T�`�W	�O[ݹ��'&LF�qϫ�i��L��x׽��M��C�9%��Ǣ��3f�pߋd��Re>B����%(ɶ�"�qW��қ�ħ}�f
 a8���{���:�\bo[|j=�ua��t'��S{rbr��-e�-"@����;�k����&]8�����E�*���j�������D=������t7Z?�R�Q���a&�)�?�e�v� �ƥ4Z����\��Ӛ�����xE�Ԕ��-��PjFJ�e���pߢ�i��S�G?r�"!S>��[msl����nc���j�t�y�����&[��c*ϟ�M��^��p�aY�>`���ŁyY��ܡL�v��%X�'����-�iE~�Dq5Q$��^�����>4�b���)\TV���g���<�tAN)\ � �a�'��ՠ�1�%�ޮ02��w¾�ٛ�V�� !�EY`O��[m���C�� r��C�{=҃�����KD��Vq�����2������V�GiNR�s�(��bݣ2����#��e�cH��۶��9;b���#����Y�WN�Nkxx5�&�	*<��-�O2.o�����t�:���A�2\��L��Wm�/�R����v�S-�}V�ƺ.��Io�i�X�J��jG���X��{C��m� �D��(����P�Ds:dnݚ���Kj�
�=Sn�.*��@sp�^MI��Y��4�*�>�L�ȊN�����	7nab��z)�/�k�2���4���$�1O��AI�YĦyv�BXLڃ�R�7r�ىd�uS�RO�����hu�����Fۋ����X�{j�rJu�+]��U6Z�m}�hA�Z%�}����m���������R�m�`W�wO	�����⽇m+1"d��\C�x3��X\�����7�R+�]虝��ԡi�a�i�=�h�����[��V��[6R�Ϗa��Vx<g��8��L�?͢�ؗ�O�� � �B�%�����ՙ^X��Ƭ>e����>}����GƔík�|�d����A�®�тÍ�x�<)�F��YX��r���	o�	���!b�+AG�k�b%�`�<��]|�
����ET�3N�m�}�}j�����ϗ��ۙ�UA�Z�|S���<H^��=^?w���Fvƴl�k�{�'@L��d�pB��`�����$	ћ�`~O:*`>��qA7!�� 4]EVԘ��7EbA�k��U��z7�P�X��O��L��6숋����B	�|���^�}^s�ǉ}��&����Bzm�xL�G'���Wy�N
�[��mD�Ƈ~h��QÃi�~?��4}NiV��o+uC�7�5��=���&b��",y~�7�� �,�W&���,;����L�_ĳ����Ch#�W���
����K�d�j��w>��Cc@�m䎈�4A;�ɿe���C-��{�e_��c7�T�h�����U"�v:�;�iY�D_|R$&�cPi���W�v���i���k��F#�X|��TWF�B���D������YZ~�p��� J�d����JA�Y�z�����`��j�F%}"u��N�` 52�\*sNL�vQ��}��(�.�3�M��d���|Iz�,�c�?��FO��͌�ʠ]}U�D�"�N(4z��+Hۭs�KL�ǡzn����yr9����H2_jq(����9�WY�)��5Y��k�
��������Ϝ�]��缬��?�&	p��#=F��U^r�0|�-�e�3�'�`�9	JK�,}BUy�<o���(��o���M�&zѩ&DyO,Ȧs�E��$N�vP|8�L@�RS�m�W4�<�A�[8�tdh��6@���%j��3�T_�Ȼ�"�����2�+�Q5m�ā�o���C ��\�*lvs�uXk�[��7$n�r���F��"<���W�m|���>/�Pmf&������TvA��y3x�r�M�N�y��Ϗ���$�~�)��n��F��X)�e���Tu��%a@4\&%�g��t6��-�&\�	�!�-=n�8O�PJ���/���g(��o�V�@Jd��/�1�I�����o� >�<�ں���B����A�%���؅ݣ!9v7��ey�JU�#���.��:Km�'��x�:���.�/n6�v�֟b��o�Csņ�p�����z��ROA�'�ȅ:]p�g#��bv?�5@�X^"g�x�-�{Z���P��&�^k	h��u��)�����my�Z�H	=(f��wC"�W_?�;ow��8���s�d��L�+�1��ͦ�����^r�eM�_�����B˰Io�9Lf��at`�kD�,#l�I�p�\�6���
��`d��5�������$�A�	֮WE��HX	~>a
$���Iٟ�uC�QJX����'�E6�5g۽�D3q���b|֓����Q��5�A�]Y�4N�n�w��KCj��,�=˂lžUB/����� ����`�k�e���M�t��x��>V��d~�(��6�_n�]C'�����H��xM�$��M��Ӧ�<(ڢ�2�40���V��ի]3Qk��ZD��D��@6��Iy��A�q"�!�<&�(u�F˘;#�g�|�Il�s��7�Ӄǩ҆��, ����/-���+ޑ�� �Ϻ$�a�M��I��k1>�lc5&,��JzS�����G�8L�e��dIVR6nn�(U"̸�*>��Q��;���ص9}�tղ@�_�%�ew9���ÃMQ-zK����aZK��3R'��߄�E��g,h�<�����W�] )-z;KR��7-�|�SX�0����Gk\��L��宊C����CWX���+�����|��N�����p+���Kī���8�Xk�'M\��X�Iu�7�K��l0�:� �����^�^w��5yG�����\��ClZ��x��1d�a)�P����p+��4	SߛKI^t�l�Ec_j���RԱ�#��la�ʇ�
�J� ~R�i4��E��p��/̈�jV�����4�c�$z9�%{��ƺ�-MʗWê��]�b�2W��
p��"�]�v�+���w����m�ð�X�Y���7�(q�A1�1,)G��D�}�c�k��Xz/W�F��95%4��� $���d�צ���w#|4���଺��|>�s>�Z�Ve�[��7q�;]4x�L�h�k4�[=HQ}5�U��ί4�}��;do����,-sbT|��x���9X�C����]]�L$���E_]5�sJ�vK۔�6��3��g��Q�����yt8����%�E��{���������8��7 ��a��U5VN���--�{1&=w~�ɐ�j�E�`��i�+�I���������$�=ɡw$�חF!z�y�
��
j)�������� �VO	����������Up���㖇�U.��a���<���s�G�'�	�P��w��AB5���JE=>����$��e� t�P�5O%�obQm=�����b�����Bu*���/���Sr�L���?ߎMn*� �c�b�4�HJ�)�w���ޤ��cD���41�m�p����BhwM�h�a�>Ȣ�T��N����J�9N<\-^��]b�K���Q�����F�pt)�� oH|�_�"��uG�2
�{�5��ӤL��!�֫��o V	�j�9R 1�M=Ҕ��o���a]cʐCב�����|\��-��eJ%�<�'qc$v2O��H�d��3"
�1�&�&����C�f�1$��pRz�z�#�Ľc5�Ė�$x5ᰝ�m?�_<����J��YQS&{�
Xo���S��B������IZ� =��co��9�,t����O�a���$�
��cΪcck���z�/,�����G�4�	ڶ,�:�1#~(���91�e���
0N<~,��..�@���Q�_&_C��~_*�0�d`#�4f�Iײ#�t���8z��?Ƅ	?>��Y�����0��wG�}|T�:;�K�!2��HؐQ �J�Q$�C�����Y@{�w9��}��</�α/��?��*�{Uܠ�Q�(~P��|����"<��)�V�}��\��9A`�Ḳ�C�-�
6�t����8�ſЇnS�U}����#�'�,����Ѕ;�f]��ivEq��)�kL����ߑ}R�)�h�|�W�t���ɨ)Q8m$DՠĴ�$f�ڋ�Z��P�ry�W�|H"J
�҂� gO���~����{A6JL�W�T>b���������x��)��oay��5��c�ϕKvǓ TpdkQt�ԛ�h��ե<�V�?�R�7p(���K>��"�'����^2\��_m���|�Z��l���}t,��k�.lp��n`�Z��j��gP�{�	v֭��N��<1�c�H��'b9�'��L~N��"'�j&�d��Vڗ:cȰ|(��1�r����<=�(�e5s����\������Ln�*�2hT8�[3�;�gn�����.a�
����(�v�ۦ��<\0�O��Nd��X	-���6l�ȕ� @����J��*;��,넞����Q'�pt�aZ;����kA>��BN�>L���h<��<���7)�r�+lp���%y=*BZ�D��Eԟ�D�m����CL�:�����Zq�I8��Ιy���Yq���z�:ǧHx7�7ʹM\m��_0�� ��M���:��c�i�#w�� bڤ>G�~�1mA���L�'�����$�:�� f��]�d:���A"LhN���|��#A%�b7Є�K[�?^ŵ�o�K�#ͨB�*#ծ��!|I:�κ���ώ�u�xI�ޤ����:������ű�Z�m@��}p:�ܬ�?���6vi㾵wz���MI��>��P#p�6Ͷ�
�����ZcK�N����W� 9���o#���(��e�����&;)M�ԣ�/>�)��d���1�9�+�C���6��?S��aF���jt�$Q8�7v�DO�V�&�[�>�A�}گP��8����F�A�Õ�
r�7YY �/rct���i��3��[�~!��~Th{�S��z�6�s>�trO�t�bO^�u�K�w[MrTkр>Ն���uwi���/J�/�"�6D&�������:0!E�o�]g�S��mLVo��&E��lxPky7b]k�w����Z���la�g��X`�;І:���B9f()d'�-S��TJ��T�Y�;P���j�1���wt��%���ѐ(�A~v�O��X��^�����<�DOH���_�G�^��?#�|�T�
#��JS���K_�i�o0��z�l�ә��QV��(7IG�CFo���E��
؜J�|����SNv[�%�:JN�I)�\�3����<wS��V>��䋤P��#�_Z1�s��[��T�����%}��􃫳w. ��E�������Ly�4n�O���+ #���j�]�ޜ�Fq|A!=NF��[Z]�8,����Jj$���V��b�!�Um�tE���\Ɋ&�B?����>���mJ֙�5��4AU�p}��=��F��)��y}��Zx'88���3�=\�����i>�w5]^�sr�{��vR]�/��Pp/�����p��!s�Ʀ,a4h`BW���P/�!�D��pNM�Ԝk\o��Vh�h��g-$B��%���{���ۓ�M�tҞ�'w6��n@��I��J�<d��g�<��\��R�8`7d�U�'��Eކ=Z�����Q<xf��Z�;C�U��6T��M�9-�Vx�)��$���K��Y�G��Ebl�ϋ��p(�]�Oc�3[50��j��[�P���[������?���(����-�G�fVL�rq�x"׷��:P@�z��I��qb�V�&7I������rO�=��qu�����w��*D0�}+��Fq������|�(�F�8H�#�k����zAN����{�\+�t�=�4^�����3C<��t�a
KD-���Kt�j誥!E�`S��ʕ\n��L�
>KXX��%�x�3����	�R����:^�2�)���B�C�"�n ��Ө��]���ib��m�x%v�ܿ;�9Z@���k�����4�F#\Su�@�D.z^�c�	W�R�=ד�X�2əs�j����z�x���Z~�>rPU�|m�����*9KO:�G0�����SG�k���g�/*��1��+?
�u�a4'�&��&Q:��������Rp�A=��i��Ѩ��]y�ZW���Γ�����q�Ӂ����PU�V9�d����a��^�AZXVV�)���|��rg���^3J�uP̒V^B�0���f�=?nׯc����g�9��#��L� ɳxy�O�N��q���ڀݩ�#�[�O�ʽ��I>s��G�Oﱛ���]`l��S���M?��^\�����v�%��}:�dφ��"h}����&�Ҙ�KU��4Ʌ���y�%A����/�3� 1��0i+��F%����y`m�ǩ&P�a�42.��$�ӻg$g��6[F�<��tnr�rR������уr�i���Q���͵�I��0�>+>y��=��Ps\�	2�ٝ:3��y�wq߄%�l���~�c�5����qq;�hx���Bai'f ���I��c�1�R�<=b2��xa`Դ�d��;a7��C�l@�6f�����t�4﬩�%T����d���a~/���Z*:찟)�fk�-����8{��e.��� ���k	2N$���
T�6��mv��hm��wu�ƨ0��Ȩ�ƕ��ŋ��|7�94�2�&�[����eܲ,�iλ��_��7,a����x�=��$�g�>��~�{ ��X%ny���t�)RC�����[X�u0Nٱ#����╰KQ�o��K�V���14x�b�����g�m4r`�?����;�BB�/F(c��X#G�Y=�I������u�l����N`�i��ǋ�V�~6b{�C��4�����'x�
ŘZ�+���.��Y�V1�tMe;B������|欪&�V��Q������G�Q~�z m�ڣ�<�8��k)�$'&j��Q=���zլgN.���w�C7��]��SxS����^3�{W���-o /�Z�ɕ���>|�`�\��Ef }�~�7��Z]���<��7j~"r����LΒ��O��H]���=0j��ٴ��$K���pʼ�x\O�
�����d��"��O�ت�b����y��'�L($���G�)�����F���l�I�nً�+��73}*AP��N$}G�ju2R6�D� �u��)��c1��ß����b��)���x��R�ʂ݉W1#}�ϡi���z"Rƒ������T�)2�g��	�Yl44�mK$���}�jc�vP%E�b
u�>���8af���كXwM�@gCh��ͨ�8�t��茊��� 
�W�rߒ
C����_HxFt9�$NX�ؿ�c�-x�<�8��A�/}nu���_U�t��-)����3�';�ߙ�S�m�PAL,b�������R���ܻ�zB��k�N�DÈ���~�#����"M'W̌��9)��/�����_72��bm'���ϫF9�j�����p�S@6,>���Z5� ��&��]�&h�R�S��tZ-��TRa��Jm�&m]��؎r7�C!�X��a���-����ᶠ���.��i�¢ofH��2,[P�ZsPʆ#�7��ٞ	���N�x�IJ��a����L:����/Qc ��o6�%.����C�6�(|��Ų����fMѭ��p��ڌ�K�(�����LH|���4U	�{q1a_�����Sט��������$Z�L^�K^۪rs�-7Ҫ����+f��<�>t��ѷ��q�3x�U����[�]o��[Kam9C+��J˒57gC�c�(�5��`@E_���f2X��`�"q즾�_��4sRVr���0u�<@�&�V��S>,.�߮��;�@��ub�H���C�J��ݖ7��/���Յ�uLwa|�Sh�msW�cs7�:�I1������1Ϭ�II~Z��<�k���u�Fӥb,k���53=_���-q3��B������0�{��tvR���³��q�O7�<�.��!c!#�X��"'y��ֳ��GC^$Z)�ү�ɾ/�*:.8���[��3��|�Up�׋��e'��Q�aqQ��Q:Q����D��-c�P;�Q��?�_<�	��Z�<`Ѓ�tQ��*���5��w�0��՜.5OT�W}>U�Ŭ�{Kz�[;�V�
[rB�7q�?i�r4j�Ҵ*�����7��v�mJ��1�_Iqn@���Ooϱa�u��Y��|'��l��Nv�^����Z�B�3�N�we(�j��g~d]�O_�GHOߖ�ugH�����[�e+o�;��ף�ǵ#^�����jg=�
�>�}-����h-�v�V�a������W7��N�lײָ����"?�Y)��}�xuU���&�	�x�$��;�[8��l����\��xq\����"n�az�{��39�?PZm��?'��¹ �E�r �O�7tFx��13�w�#�?Tb�=^�z69���vdi����L�('�D���}���:'_��l�s&����&�Lx@r%2��o:�� v��ڤ�|��]�"����|�X��A�� ��[���y���1�����W6��[��ܕ@(�%��D�<���pK�(#� IjO��j˄�8^3��K2����R\ 0����pX��,1$Ȩ�)ܴ��=�d.��<���v�ٟ�l������I	�ɕ�;X@�`1���M����0���<VxRn��q�^����ʽP��	��$�$@R>
�ڔ�hSg^�la.s��?FA�����l�q�T���k[���p�3�j�h^p��������M4v�0�6�x.��vd��fE,�`mWnk:���}*��*(�mF(l +"��5U�0��J��m��Ot"b�wR��^'R�j���)��gL��`)a��3�����@��I�)s@���Z�օ�`b	������)9��~n6zɥ�|P�U��yQ�3�&?�P�X��Ax��B��p+����5��`�F��g��.��q	=�u��B�Պ�~���p���z�qg��a�Q9�^�SY;���v���b���]�W�8���_I���x�gڋ�%g5�-E����w��t�'S��wm��hhׂ��W��i+I�V���^� �e�p_�a�+r�垲�X�>�RI�j��Y^\�B��Y��"o|4t�&�+�@����&��8������Q�`77�mX�D{H�ta���?�}D�q�sb&~�o�3}�R=�]ޅ	�@\�ڣ%ٳuXaCW1�<?��k 9.�`�(rpU���|c=�8�=�����O.��	�+yzcT-�1EvʶJm�cW]W������<Z-[˃^\�w��>�)y�^���H�.C����ַc	�4s7��v��cu�%3�
H}�WP�m1O����I_�����:����J-W���������+����!nB{-k������S.����r�����q�A;��C����$�6�_���m�hu 3L5��	8��=�\ٻ٩��$����b�G�?���-�#c�<��z��o�ݳ|6	)��E?Lr�A��&����5��>lMq�r ~\�e��\wPF��یe5�Nz��������%�D�8)%5Z8��b������|�=�Mt��1��c�����ۖ�DT���8�����<���.��I���Z����^@�m��FIV&*H_Ly�m���+��Aw� �!]Scs����|9&��-:iZO�O)���3me�iTa��m�H�1nw� :�[�8-��`�Ʉ��/�
cX�#e�OFsbC����NmL.~ s�V�[G)����΢�&sGQ��9��w�+"G�[��N!C�~.6����W��_��M)2��:-A8Q�uc�@��qF�}X���,�׼��R����,��u),���hJ�D(>ȧ�|�zs�|��8:�>�k�㫌�G�?p���n.�ʅ���_�;�s2��gO�?��F�'99'#hUC��Q��=���*�ȁ�_�J؁U�{ep|�D��H@x��m?}P.$��r5oK=*�PjB{�j����z7f�>F���{b����f��I��LD<�j�m�?;��I��{�B��ԋ+��c��EC�����1�����3P֭|,X�#��&�Olj^�1+�ƁZkV%tO�W��.��lq�˅2�����	/����R�!�B�������+=�6�\�W��
��=�\n�Qҝ����4&�������|����e�^�'r�o��ժ۳����o,�n\����o�6֏�o1.�e0�e�ޡ�cvHA��C��7h����3R���ߔ�O�N�#x=��>�f�
=-�HT\�0'���Eع-/u��o7��/M!��>���}�4���J���v>�Fe��B��=Hlx�s�PU����&n����/�Rީ.R��"���N��2���ZՀ�
͜��A�8^Ix=�~K� ��Ŷ����6��m�j:��t����菅�(Fv	G�(�C�:�c��!#���U���޳ʞ n%�x��LN�X�ϼ�Nd����'��),�"H��`�D��BN�FA^]�V@E�S��W�g��q"#�a��QI$Z���]�tn����$��2.ȧ�������߯��!��qn0��#�����䀹���Y��8BZ���Ԃ�Cy�p�����vm�Z���q*B�+8�����_l�z�pp��B���a��]߾ʧ'{b{��.�<���sL�p��vX=Ӆ��"��$�2b���!y��	؝�k&w=䦥�Z�Q��t�o��E�3����>(hy�4D���
86K9
���1ic��#0�-�2O������ۍΰl�#i�#\n�L F2:)�*�$,�2s���w��N�� kX�[$����*����%��+L�ȉ��6ތ�do�J?5%⎪ڣ1=���b	��)Y�MA�8<���󳷓���;�UK3���p��j�����ǜv�ת����5��7����Bi(_��ګ$.��,d��ag�g�xl �[�\�o	l@R8�	��J�Cƒ�R���v8e��yId h��&9Y�K�5V�:m4���SH��I}l@�x �s%�H�z53�h�Aܮ�������e����,.�^�Ƴ�Z�ىs�B.��WsԘ^�>"�m�Y}~��/]���UB���E�`���d�wMe*f�e%`�:~/�q����-_�AVl��l�	�ۛf�1��)��L9�����9���U]�0�q^���̕��ݞ�[3P`�t��x�?(�x��2�%C���8��6*3(Rw�)ci�~�"�"J�K6�0�/�1D�4~ӣM����l�()�i�4"x�WS��t~B܎=����)i�	Aȹ��s�@�b�X�@�5�3V3�`���w\m���
Rϰ9$�h �c��]���})�_s4�0������L�9i�B��CMC-EQy���2'�`S�'���a�O������J�S�/��)� �}&P���o�u@�Ѯ�X<xz�,�	b���K�Qh�ǧ�!hnjgFN�|e���q��Fz�V�����jU�Bm�L���������c�~��-ψ��o��
��DW������`��F3���e�>:������Uf;L��� B ّ� 
�m�r��f�4E�� �vrk�Թ[��X~�hȖ�-��.���mB�Ǫ���S0�|���%z�mVd�f��\���]ivb''����CO����$�Ȭ��ZQC��EL_�2 ��@)���K�p�I-H;���NX�\xJ>�6،Q��^�w&��dŌ��M��x9�T1����5*;'5��0�sV���݊n+����Bg�ꆹg��O�7'�$p��i����-�?T!���8��t�sT ~X�,��-&Á�d��)�ų$��+�!�2��d�4�(K�qB�:Z�h��`��Cl�8W'�����b���*f��
�D	1�i����7e�Ԥ��y�b��ӫ}*R���S��ag�]��V��}o�j;���so@{��*l�`X.����:���{�x���V�W2�l��j��K����<�>C,�a"Lg^�K��f0�6K��6��i�������A'{�.G@ ڳ��}�-����>�����E��9?ȇ�x�4�
��)�*}?~GYd乓��6� |rj����1�k�P�z_T^��h���\CM��%��ښ��- ��r��b3Jmݝ,>]7�^(E(���d���;�T'~�%5�X|����a����ɮ�X� |���s�]n��
�м��հ�S����Er��W�B�\����c0 ��Q���(�F�h��?��^����CؒYxƝXz[ʊ.�J�|��T�K4W-�Y躞���$&�T�Pڅ<��cs��v1��3��>li*�8�޺]���t�E)��x��BiS���:��8u��*u=�tZ��󆀊���t6��ہ���~N��mO���)(-j2-Cg%����݅����i9J����œ�W+�!?*�"�����iä���mdH�H��s�jZ'�x���*�~�ju�`���i*��|�63��_�.���e!�ZF+1=��g�c�y�j� g/)��i3
��yd�e��*�Dʍ�F������'��.�T�S�we�1ԡ��:t�X��t9�3p��& y7��^5��V͇֘�#"�4��6�Y7mX��,�VM �%��eeY�*����aIx��	MH;��~���텘kc�Eo=?VӨ/�{ѥZ}�����V�<#��Q����!�5+���^dL�Q�;��lQ��bM�du���v6	&&,�0WTM[N<" 6|�n���}�[��s29z^��JJy���ڢ`R��]j*8�s �h:ְ�l%���'~��nE��$���\�3��z�&k�>U0��ڭ�CV|~���X䧊���n�i��� k ���G*M3����G���`�UI��;����fk��aآ��`-Xc�U�
���(��l&�5���e�2��3�QKb�M7�x�Č�����\b��������	r<[��9N�'�-���w�{���p��%Z��k"�����F:��ժ (q�
+��ܿ����\�XC��轙�*K�cӒX�u�&(s�<�܃̝�d�.�Uhc�\�1@G'3��*��TF"�K����G�F�j�љ�+�Zx���uS�p<Ĭ�\�O����|��3�ؼ8A��9��*Q�Nީ���DC�e����3O�4��G��Y����f,���N�6����t<!hsҳR̮��かpa�U ���'>�4Ak�����?�~^\�@��8,aY~[�b�㍓jNٿ�����gͪw.G��I��s5X6�y��l��G͍�WER�	V�?�f��ـuGD6Q��D��Y�-`��L�E � �n躵+@��Q��mZ�=�����զ�q4F�G�aNI ��м��R#V��P��hW��(����N���r$�6p��(�j�i����A�(p�`�3��k�d�;P���㚍a���/�do?��V�/ׅ�;����5[�s��p��~]x�=����Y���S�3���xt�K"��u�k}=�4$��O}��R��Αz�A$�\@�%���fi�j�;X(Ԕ2�6s8T^�j�8�kq]��|-����$9���=7��JO��T��@f�dV�xnG��TL�P�1������4����Q{���GI��޺��po�� ��W"V�n�^���ϐvs����B�Z�ϕ�t;&���ؼ�|dj��E�6��T$�,�&��U1�q�Bk�g։��e*�ȣ��'cg�����G0_��[�=�QN=2����_�ic�w&+T��rc݅�����k����or�_�J���Zl�	7:����M�,V��5�r�w�v��SrM���^[���a���E�����}��Ƶ����̯q����L��IE:�G�9���IY����y�� jNv�l��d����*F�z|��>�C�qJ��Hoq�yU]CC�-��G���|M����Fƍg�d��p�'�vgp�×V).�N9N2�
��;q`zc��Mn�-�y�aP�v��	���4�e>�p7 ����{�ȳ������%��8�Trr������v|$�C#BK6��a��~��T���e�o�:H��M���o�'q��k ��/�?�hj)�L98R�m�}����(�7�������x���`bVB쵟�g��5Xbǟ��`��Cd�py���mr��9�`vB���՞c�=cp��� @��VF̐�e"��� 8�Z�Е��e�'+�^	��}�cz� L������h��d˳/n��V��9�t��[��)?VG�
A���={�Ü��,rە�D��Hk�5��ZY$�ί�\��d���]�I�U�L{"Z̴��Tz�x�<_��\�5(WRs��
�<�:j=��Tu��.�7D*�tNj,�i�o�C��=�m���fr���kK��]�ө��7fc��N�4V۩��[��=�_�|Ʀ�-�l���x��	Њ���c�˞O�j!�|\�������:T�7�g������;��� 4�[��lG\�a�|�Fg'bvg��ab���@C��*��	��t�M��ɻ.U!�,o)C��c|b#��ri�h�\_����Qл��Y�+}E�0ȟD������5�e�5}�W����1��0��B��ȅ?/�MC����*}@���y�%�m������Czp:s2����="��7ة�XI�U��(���]G/��Y6�_ͭ�7n= �1��a#�ɦ��:�9N#�I�`98�u�7��>~���.���G��up�K���̬�`)�_��6�G
N31����R�^�1��+���E	�6�7�S!�w�z�?��[�~�򯪻�}�K鱯�
\�7�v�� F]J����:�a9/p�r��Z�%<�
�x ��=�@�6�t�QZ�O�[��^Q�kӡZ�E��>u��`�(�z+˚?����G�9��`n�2�&2㆝�c�Lu�< 5��N�U~O��f�L�r���H쐊,�]��5H#��6'����6k�����aJ�>4z�~ZFEY@H����C���3���e���	}g�N�;����櫳�2��!'��%ľt�	4:��d����=���5rϠN�����k28�Rr|�&l?�{�.p��ka؇�������0Z����	ן���&8MR({Zk#Vh����D����O>��B!Ƕ�d��q���pʇY�c( #���KW��s��sX�u{c�X���܈ѽ�?
��gQ5oͅ�m�|^4�b�}@\�v|H�W���}P�X�hY|[Ě�ْ�*w�щ,$��M��M$��Q�?h�B�|����Jd5������dzUZM�ԇU ���I�KOZ����2xmT����E|ȟDƬ	�{Հ���BK�� v�N���Hv��,X0�N�������KdS����ȵ�"��ƴ0�����#9��*z��G��fτY��.��=6��bh!�~Q�5q��ޓi��~�`6&�E�+����uݰ9���څ�3O�S��h2�N\�}
� 0  ����s�`T|��{�Y���\��vL��}�Z67|Ȣ)#�As�?:����ل׮�&qz�w�������|ÿ}}~���v��������S6}��|�W��n
H��K�	��5�#�E$�6;s�}���я
�=�!F]o,�������48�C�"��;Na� O���9�(�Sj{șY �3��_'e­��r�'v����]}�}X=Z*���핍��S>�V6����c�i����?��p�T����Ps���&�@�](_�����8_>�,���꼘��O�Qs����خ�&�����!=�
����!�d���5iT��3�����/��_a!�1�޽�j�έ����0�&/�鿶��M���u���5B�˙}Ե�Y>p;�l��﫜�+�'מ}/�M�	Nj�R �a�b�j�,���#�R�f���V�5F�*�I���
�ѵ���l	!(��[c�{�D�<$�u]\�"�N����|R,��U	~�l��=Zj~�� =+��R˼/˿���wp��,�$���e{dh<���%R����Dy��a�n�'�z���I�����R@UYb}n���<�̴H��T=fi"��`�1��P��6J�ta�R���$S���k`T�k��z�}����_)8�+�J���D'���UdH��ܐ�6�$���Mʹ$�/�틠�һ�f`XaHI�5ZN$�NP��w[��	(����q�����d!h���lT�Ї������脣��!�|Yb�r*�M����k��։�hj�����4��`Fp�@�m~>qb0�R��Z>.Mj'	!)̚��� ��*�T�ɰT�Y^6nK�>�u�
�B����<��υ�{��eZ�k4�aHH��չ?���4��|(:�@D��G�8V�f1����]�o)��Pz�r�k�����r��u�D*7����H�5C�܇��栳5*��@t$&{jS��"v\�9_ص�ErP��GʾO�o��ؒ
�W>�n��\�K�9��.�L�NDKa�m�8�L�2���5�q��Y�]�*�b�S/�[�t)rR��ٹE � ;���р�^r01ŃPa��ߏ��Y�NL�T��;�(��A�,"�� ��i3���h�6*1�XN9�k����C�Z��I,[=$���MڿT~G(�9�*��Y�o��U��)�sV@y�3�:=�R/����&�<�Gk`�K�6u�~W��{>�u����W������j�w�k����:")7p�6TxH���n�I��|v�E��&0�>��*�p<�����$K����{lx����Nĝ�3�������{�F�iE��8)�4@��3q����Ror`�� +��pGJi��7yEA,��ۯ�#;ȝ8���^�� ��X�e��D�%��Ǿ� �.���V�a�R���>V�Q:f��v(E����RM�X�w�g,��B%�M)C 8�0S�\3�C�|���	C��Ч�[�w�	8��U*8���ֳ����*�q�Zxw��]^e�9�y�/.f��&� �&+-a��0��d�9#�Mْ��q��+g�ϸk��mr�����

�Z����Ҍ����޾�G�w�d?Ț�K߁��V������˧��Ceϔ�&�<3oc;l*|��p
�\�9�o0ˀD?&C�J�E��U,��C��� $�&�)�����1	I��Y�� �_���I���e9�c^�$ƭ�~z�B��X9�k(�+��ݩ�X ���_��D�,E10��>�����d��[������s�ND+�y�����ޓe
&%04j��X~�?򌓉שg�CUk([��zN]��*c�(3PY�a�9r��Tڴ��v���2� ��bBy2y-����8�-�pk�F�0���Uy��Qv�i�Ї��$�j'��_�XO���)��T}��V8�t�+���ĶHՀ0������Ӗ�|H�9rT��݁ר@� �O�=���!�=���_x}�k8��^�FV�-&�;�r��Y��+A�H��I�?��~�!�ҹ�G蚲X�YL u����@���| �����p{If癒-����.�
c��'��e}y�x�^6��7��jC��֒%�;���1e�TH���c��e�C�0���]]TGF�#��4�u��On�V,Ђ��[��� �2���Q�~$s������+�ü1�i*e�'ĳ�	�@3��"Q�Z���GW �\2���#0h<t��ܶ�G�8m�@h������|�P���*�/��
�4��%�� #���j!���!�[t��9��:��I_�	\�(p<*�C=��7Q�\XU�P�e(bm���\J�5d��5��I��tA`��w����93�o�Hn��:��1Ɛ�WӢ��Qz����b(�b~-}j��AC�f�]�Z�?�lѲ�|�0�=�%9���)��=� �^�P2".M���g�՗�_�Z��$�o�������Ɖ �W_�KF���� ����(�b����(t6�VA�����4�*L;�yҟ{�� �N��6lp3���JM�S�aH`[ ��J�!�m'�f��U] �5�S���e�T���ΣZ`LY�qJ�f ]S<x�������GJ�_8�����l������$wֆz�V�aYާ%�����Jp�%(�#�R���Kf ���O�����[��û�Ma�	���C�L�7��(��+L����s-9�z�KԆ�(A�~���p�_��mKPO�CA<�l!�h�P�
�q���z~��Y!��>�V1���J7�7	����p�#O�!����
eQ�kJQ?E��Mh�S�L
pP�.d�W��j�Ǖ���9:٤���U�4�(
�����y27��Ǉ޾JZ���[����J��i;͖L�l��c�U�Q�S7'Xy ����f��cҖ-�c��Ν�ѕ�Ȏ�%�s�n�}g[�֜�ш�ů��"V
� �uH� �r�IQ��wu�+���E�0�9K^�w��(,"���&��%;x�WH����\$��0 CX��ʐ�������oZCM���tȬ�vh$q-(��݋�L�8���	�*]��=��{���̢8"bL���Sn��7CS'�	&��1&U�,";bHf�4�+�(
:2�`�ֺ���O��#�eW �����L�I'��12e�4�4��O�1b#-�N�hA6uV��Z�/_�];I�ү��M׵j�M�C�,,`%���<������qxw���d����D��iyۛh�O婏;�nq�(؝t���;�e��1L�m
��Yt~%���*�̙$��&��*7	Yd\�F��ӟ��lƭ�G��	���;	>MK5�a�%�+E�M�
R�k����|�u�f=t#�h��`�o�J����ߦV���H�#�Q����c��~X����0�caz^�㢟x�ͼ��pgm��A�Sz��Q)�n$�:��}	i��WgE��p$n�"�d:������}5�hYlҽ4��_��7>ꉣ���2F�\�����>IZ�2�	���$����-��O��dʕ{�9�"����(U��@hN��w��ܒ�V6��$�3����u�H���y�CZ����bWÿ����ި.��>g��z�8��e�Cc��m*�h��N+���u��m��.�y��CA��E�e`�@�K�w!�^|y=PN��k�rQ�^���/�]r��ZD��nX ����6��c���W�:ϱ�$7Z��J� �^|"Y̮�]`�:�0�e��f�HEd��	�A+J���uX����~H�A(�;�1�k�~5�MY�X|M��?�t9?�_+^������k����x�*9%��v;"�c��P���Ikz�#���t���E��[��������F��P?n�zS��=���% ��lS	��������ˉ}�O��잔� S���`ּ{1�ć��қY�ә����b�=���a� ���� �r<M��a��e��E���G�x��D<I׼��I�c��-��^Rnb�+�CՖ��+ru��ȃ� �} ���=��Ś���Dz4"�>½��/w�ct#�z��*}�BIy�G~�����8�w3�G���;���gm�"-µԥ˖5�xaW����D����5�����\����=2F̞�\J��ȫ)���`���,"+t���{����.N;e����*5:4+�A-T4˦_z�t���F�J���M2X���a;{�M�����C�/Ǫ����� �63�%0>g]�v��ڧEK�ƾ|��'%�����C�S�k�Tc0d��Ы�Z#���{Źֿ|��ް��g�\����R��;��c��tF@��-l|	�I'�-��H��jΪ.Eu@�<BD����*}�\:���*��(�6M/C�7c�,s���(�l;
��n�٩#�j������ ������,�g4�_�����{E�X�����$m?��KJ{�!����eShD��B�ݽ(��-�1l�8dE�����NdV��=�~5�V��	0���/=%�{1�[=孙޲DB�}r�g�͇�����0�Q��rY1�Q+Q�%'`D�ۀ�x�VS����'8��;��˒�����*�;I��d��n,`���c}��m�]բ�6��=Y�����sL�ǟ�C{��:c2�q�>X�o�^l�Ee����N��+�s�p�.&�>CS���bY"P��WS��3�ko�*�|,��v�d�Y�v$T��i+��3�k:l��9C���k���y27�s^�� ���h�S��A���Nݮ����~���ú�c��=Į���Z�N+����H��"U� A�/�	2������?2�ާ_Z&	��NT4Q�d��>��<��@�v�o6V	:D�Z��v\�e���y޽��\JK����W�u#�RfK��A���^^�/]��Mַ��{�q�.��P�Ȅa3P��I���^��k?Gm9�2�"�;S��sՓT���%��9`�����.��\I�	�����c�m�ԑ�X�G!,�ϡ��0βŏP�q��+{/�z�u�Us)�(h9x O��� +1��$��v�R*��'=Ug����TsV��ز{��o& ��@��M�E�('4f�ˑ=���b
�dg�s<j���a�@!�� T���m�ɺ3�ĜKj{��> �O��Ի�cՖx'=�TG�0`+.q����iP:�c*)��Bc����>��Ĕ�>9��1��̵E�ը�^�����I�*a���-9=M=*ґ������}lb�v*��, +�{�f�cU�
�O^�CO���j�Jw�})<3�rJWtUH�Q���
�[hO��wEg���=G]1p�Gł��͈W��ۏ�1�����K��k��$��90�$L+�Qs�E5���ь���e%	���Z��ؼ.�Uj-AkX���q�@P5�c��U��I�;G!������5�#�M��U,uz�zH�Gf�JA�	B��{g,�'��}D^$w� �j/$YF]�=��O�*��_���"V�^�S�C�_����Y�����LV_��U�*��З�v�����I�	)� �&m�o� hn�7ly��m>
6�KD9�2HI�5�Q�8�R����e��;���.��N�'Ǹ�J������iL>�����U��ҷ�[ڟkF���H��#ϱ�U'�����6U��˻�6c�ӛ���������e�HS.݄�b���p��g`�7G��L[��j]�c�m+����d�~��5�?s�EW�D�ZҦ���c�!e��fY�71���`�ɼ��a��J�?��AL��.j��)�c�TApϘ�l&��E�e���Џ<.��`�h�JbZN�R�U���*k�ŗK�|�0COS�v�(�����YE��:$������a�/O���v�s]�f�m�[E2����.p�I!u"Nۊ�x4UB�6�%E�7jB���J�I~ĝڟ��r)t����8n&�iNu��3uɬ����^��/8�Y:���]|��-�0���O?tD�+�V��uwm�(	ٻ�;ޒ��5�g뺸��i�z�i!���޾+w��4�Hn��v=��<T��m�щ��Y�G����&c-��)^F��I�_	�}A��Jp6a˹�����B�|��ۧ�qb�!=���� �36�%�/lf��������f��}r�ZZ���C22�IVw�26.�5��c���E���_�o*S���2���:w���]�gl�N�k�4�lx�&�I�0�L�;�%$P&���]p8[0s8^�E��m�ª�c��N����Xw���Tz� JT�5c`��H��󴀬>������-�����C�]���W;M!��<���|h�B��c���+����X1����X�(J�nB_p9�sr�dY~P�
@�XᎻ��w�8K��K9������{2�){v"��p���@4*�,q·�	u�,gu#k�Jk�[���;j5�C˦�\��z�;iR�R c�?R��G����QG:���ч��3K��?('�,���ni����\����&���&`j����I��Qk%DÍ�?�U&�#ْ�8������F֐Y���cZ�i�`Un\Q[�mV+�'j�|$[�A��m�UՊn���s	~��r�շ�;�U��LM�%��s;���]��Y��*4!oF�`T� ��n�-c:��O�E��S���g��8�7�C.�b�S�4n����_�Q�ny���{3V����M?��%�lH��O]���t�Ǎ�����~r�g�GЅ�Eh�(�BJ#/'fbK�k�<�1^���f~g�ݠ�uuY'���e���\7��ݒ�tO��Ƌ���x�G�d�z�X�(ҫhs�՜nS�W���q���d�@E�\7`*y���Y~B����i�Hƍau2dZ���J���2m�S_Iv�W�.�ڰ��K�/2�i�� ×���TV�Y ��0�Dm��Zgz#}AK��]��
U�"�+��"�U��Ԟ3�1�ٌt�XJ��Dv�r���HD��~[`��A+�����T>����?��zArS�oV԰j�+������]-�>���؊@߱��:�R���G,���_��h���� ��]V�<���I�C�X�/�#U��z�nA�c��J;2.��&w!�o�XK��v�㈜�&a\Z�`tE�z�6�b�,M ��� ���4R[�ΦI���v�����Y������ɦ�Yr�a�������;zF-��GWu���:H0�+�p�O�!���7��@�[4I͹R܏8�C���>����_W
��MR��K�&��R�r�m1�_-s2�}�a�L72)X����Ԟ��R�LM2�U��to'P�i�n��n
r��B�sA�iv�?g��3B��[�/��̤�6��֠pXn��N��$k�E�P����S��8nh��Ҽ���Zd�����8��������
.ێ7b�mM��hS�B��>�ˁ,���W��/C��\p����	����%�1�����	�^�����^�q���kn(�Y�Q0O����-�h$kར?��:M�*���	!���Y�	v�L
����|w��6��E��r��4Iw�.����,���fk�dV�	ӏAiL�~iKd��uT�P&)�|{a�wy��Z��i`s��S�x��}��,�"�2�_s�l$������i�,�ʾ����uD�K��(|�G��2���;7��1��Rr���8��M);��\��R�+�0�Z�h�47�^	I��y� F`��O����\�\v�2|�T=>���Ҧ��Ź��m������������S��t��F�S�0��虘$��-�ÿ�}f��B�4O�����)��I����Ba=y���%�Th�,OA�ǀe
y��$�+䤋>�I_���w"cܧ�c8) ��(�(���A��2lܟ�>�V�)���!b��A?i�$M3��}�ȇ�*o�~\�%��.��<��Hk��ͦ$��*��xy�V;��B��S%����XH]mrRTj�����u;5�7w�'y�*P=�\��`H1�P�E`(�����B�����q�qGv�0��.�?ڼ;:��������͠Y(�*C�� Ԕs���k�Z�u�'Lv"�d�}���=0 m7^.�����x��m`ſt��uM�M�
<�����#D�@�Nn���]�
��2]J�ve�F!`�.�&����.���Ó K����L�LYE�5�䀒�{�_�S0.��z#������I{�ӌ���("+�9ˁ�Y�)�ӹ�S��c5�S�^��X�@�s�����a�V��݂�qm�6�G��5��f�w���3��3�:)�zb��c���������"�9[C!�q������nM��.�FSrX�AK�;�1�\
�Y$:����>>__��Q������&j�D��I�RO��n�[/��(��m��E��ei��8��e����9���J� #5���::ga"���A7Q�����D#|�h�ۦ��YE:���
���Ξ^u��^�O�|l� ݅��se�s�d��a�}N�TI���j�1�a�쎐�5�����@�X����6)���1l���K��j�ʌ!4۷Ix��D���Q�x-�{��L�5k���*Y�$Q�a�vD�,�t|��Qz�PrXR	|�Ȣ�K�v���'��"�,��yA�1F=�hV%0��m��3&�9k��D�-D�U�)XH�)�����(�٩j��~�e'�ᛓ$�9���(S���U���O��A��!�<Tl�tk��/$�)c��MX�}r����rË��Uzٲ���ۣY�]�ɹ��W�5�˺�f"��O]��+�%��r�$nW{�J�a$���Y��v:�����H�z���0S`�Ń�D& d"y�����!��W�ޘ�{,���E��p;��CK�.C�"�6"����^�?@�
F�Үo]g������~�F��VWФ�O\j5f
¶���s	"�D��F�����E�ars^C ֵæ��#�4��oB\"�Z9ܩ�z\/�����糓��ßc�r�����0���5�� �W�GH��`)��hz_�u�w�E���Y��S�47���	AG���,��u�B;J~��`�H%�? �5JBA�ٹb�g��� "���q
�0_&����D�u�kM%W�	ŏ�������eW$�%G�-����"�$�M_g�H�'ؚGVB�C�����xVx�{iy�����o`�̻��Deu�c��#u,������X��@��m����$�#_s|1�[, ;��>�b�cQ�W	��p �x�;���z<�/�xI�"(f�X�
�U�#"��&���rC�wl�<Dx������[D2����(�f���s��9\H���AF��S2Ga>��8��՗Ia:�bE
�>�X�*r�_��)sVo��� Q��w�_B��ۆ-O;l�18�Ƚ[i�^��$�n�N��,�r�n7�����k,��s�� �J���k9��Z�#��u��9��4]m�h!G9�.��E���#b#�ɞ}[���.�X{ '��I�z(����,NC=��Y���u1�;������w�ޜAW+���#SRo�{x~�6q_�%��jD�wi(�%��x}��]V�V��b�s��a�%&��TT��%���:��e�V)��J��?E��{�,-�Bל/��ӗ�*=���6ι^ד�D/͎�kۖ�9�y�xr?'4Q�cZ�F5]�� �»F���+Qٍ���KBRS����̡���`�5d�s9ځ��ѽ�nm��/�kΧ^S�'g'NC�T:~Na���~B�<���z�C�HDy�Wxwh[5��Fӓ4�'���i�����@D/#K����UCu�)�+��㦠$T��.J*&�~�O���1n NpBG�KD/y��1�2:1b㉲�@���\�4�A�q~�09�=`G7*�ﵵG
Ѓ����`�Y�^9K<p�8B	�N|��i��(ʘ���yF
��6Ă����+�	�e3���\�!���ߣ��$غ�+��M�c$�A�9Q<j� �;ޥ��:(h���q�k��e�݃�v�)��H���@��_Wx�֘SG_�6.8<�캠��q�cna�MB&�X�X��ͩ�*.���Z�lߎ�s�v4o�V9G
~�r�����霼�K҇�9��ߏy�}(�a�*}[~CU���kO T#Kv>(["Z�,�q�I��:��+%1��u���h���#�֙�����+uk.w���e��u*Ɛ-��M_�����}����[p��k�#�� |�&&��>��j3:Ii�`�e�Z��.:��53}���݆�hc��e�7�v�,$��ļj>��X���\Ef����[b�u?���62�nޙ��K�~�& ��{��SU��6�/N�FR��;�bp�l��L[pL�#�[��"[�[u��D�AZc��M��rs�	�f) r�>ίp=��D�O���M���7�t����;�Uc�׽��h�X5�L#�k/�U���
�����R���S��3���~��ĎU\%LM�)m�A���9�>*�2�	4�^M]�f*ގL�1������R���MYw'����=Q�3��Սxd���U��R�yo���?]��rt�����}���O�� ��sf���J�m͕�t�)J�0�m�k7��Yan��a�1���-��0�KI�=�O�H���N��{��M/��z���LE�(]��i�Z!i��7�����#��2�=l��m�W�,�"�	�U�BQﴞƞ5$8���D��-��ȲMk���2�g���ŏ8l��g����:y��,F߰�5&�3�2���п��}�s�?�(:)�~*�7|A�O'xc͘\���c��QP�� ��V�(�����x�u���V�(�0{`������=�R�<#��j�����5��q�3�s�UY��i��1~�b&G�ޏ���T*�&!�Dk����
B����\�"f14��C �;0���Ѹf7>��u)G�Bo��FFf��t$?9�0侀��̱t��J������a���v )�d��3뿕��$��|�E�C�L]�7j�ȿrp����O{C��<��ӷ����"��=�z1����B��2����]�y���%��h��	�{�}��S��w�!��G�������'�]:;��K��+�F��P�Czv��'�Acz�y	k�h�6�B�0}�_�1,;W�k��Ӑ�\�H�of>��^CcD�E
o��V�۲�|�����_0���j��-t�h"��j�t��^2�l����E��d�pVx��Ħ/Ϧ�qt��0����*�t��;��/��'?�m{`�"y��6���6�jgO'�A�&0kyM��4�.<�������<ă��i>�S�����ʸxL�D�>8�
?y��javA��ف�Ǡ"W8���t�s &��8iWƔ�8:��=���N��_�|&Dy�$�"r��/.��&���cF��?c��iI�$!� T5�Z�IB�O��"刄�' ! �c��n�^HuUV���Tk7:o�,�NUK6��P�é��NhYV��m�,U��8Zy�G$�PvV���S�m����ɸ7�:�Қ<c�'46�{\F0G�ha���_ޮ�1�����s4UP�YV���7jw��/|@WW�e����yp0J�mJ�7���"�����xS�;N����*����.��H\�@��J5V;K͊��qt�v���O�T�7�u0/w��A�k�[�Dqe����LvE�����
�.��^Rd������4�3�q"�7kc�JN*��3�+��- ���ʞۨ�E7��JPeM�`@ψ�A����c�PG��l���O��ʥe�}j���X���1נ�����i��uz�YQ������'��v�Nv�*��+�"Lc���8W����#������e��� zh�gfy��:�f�M��<���|<�d��FG���]��Eb�J
	fw����w�69��o��\�!��ls��o��P^X@��8ڇ[�k��B���?Pym�S%3���?.,����I�1�w�yɤ|�ت�,����m�Ӳ�Z��Fj��\���������É���gU�{��o�'y��f��țg�`�;�_��(!&�H��N�1%:5�#��qFݸ�}�x���{��P��g�=m��
,�ػ�
z̡���A�_U�r��1�E/+Pr�7�\-Ŋ�X�Nצ(_�����C+��/A�]o��*˅��*s��"Bh¶4�w���B�:�G1��'�oz����e*�#��8cj����u�F���������7���@�Q(� �U�0?C�=���!��#�X�{� �d,Օ�^��b�F��U5�_ �Z�y��oc;�W:(��g>�$��x���3^8�duǱ�kE^�
��AɈ��B˶�͟SKH^���,��%Bю۱ه�!�]Wf��@m�$N�6w$�lo�ɂ���g~3g�_��ms�L���ڣp�����-��D}@�z��=��{�n��.n#��Ϫ}��?�m����`�!uA�@,�|� �~�+�4�;��nMKg0w
������<���XZ��|p4��L�!�@r����,�15^\T��ha��?b�ŵ{�s�0��tp䢦��n�<���3�{�B�i\d���u�gRoU�GyTv���b��9��Duo�xr�S�2��X �@]�o,	;���L٦4�LĲ��G�W��S����vjV�!��Rt=�JЇ��ɗҠP<�<{j����HOK��k	-���C�����ѫ����8���U�n���F:�<�3c��9e4��<�Np�4����7)$�2@˾�
3��	=;�R��,����+Ǝ����ǐG�?��j�����s~�P0����A=850^|*�i������E"�s��*�>��;5g�m�iosr�����C])���tҌE%�6�ė���#�i�[q�1�{G&EX�Y���"=�2�q�\W�G{򼍹�����giE�e���>�I��\.��ox<���O�B�a|���+��!Tܬ�Bgw�)�q���g��i�F)6g�P%�{rB�����ށ�J(<>�"�`7A4�,n���	�L7:�
�=�oN2!u���W<���28�7 ��~�vM���6���Dӆ����bi��`�W�6~�����>"��� a����6jwc^��Q����1 w8����N�����M���d��}��!�����h��ᵁ�Eg93��k���Ȱ>"�]Y�,�ϭM�Z�2�kU� �)�*a�H	�����n�O�Gmi�����r��i����N�� �7_�Y�qo5t<�)l�>��զ���(�y�Z��F�ñ�(s��C}B��L��c����V�hF*��� ;[C�7rBk<��R�Tr����[��H�xٰ�P:�څ�)ёPc�.�̯.�,A��B8x�!���L�0#��?�K�u�o�=����:;~�0�,*cw�3�|�Z[B(%��Z'�Zp�؍ZU˘hsc�U��ِg�FR����Pc-
�A��"рb�A���c�V��x��U�[�������&2�(#�Z]�i�^R�H\ͤ�H�O�>���7<]��!��SN|
 �ײSaP�����<�9���fC�'�����_�����'k��P�G٪}D[�*PY6��4%Jh�ֆ�ːL�Y�FX ٻ�3Y��z�^Nyl�����J�TSi������w�vO���X�x���Ajo��Q�,�fpwx-�GR&uͬ������ɉ���()a y�)��u�n�-q������.�xJ݋�gd���3؋*-[����;M�YϬ��j���c�n�M����������?�9AT�_$c�2�����g��h�,�I�]�*�G�M
��(�V(�]>7?����c� }-�9�A,��Q����E��y��H�S�Jj� ���٤;~?59��B8�J�"7�Bԇ ,�5��Mψ���� ڲ��#.XT`� '�-��W#A��cؼ��&a�*�K�^�4~o[wu��9������S���i0��s�J�a�;B/���X�Q긼J̞ ���`�3V[N��-r��2X�kDߟ�e��dqT�&Y6�Y��XhI�T8T��oƲ�b�T��3�|t!�-_�gNL�;���b��,V}�~W=x�5���/��d6�`e�b�s��$z?:�+�ìZZ��'=�6zF҂�K/ŝ�*�dk4���"����y�h||�nH8��J�h;䟷ҍ봪&��FfX����V��c$-޵aY��Y�5������C���\�)j �-e�YH��C��tcMY��̡0���m82�Z欁<O;�>5QV������v/��s�����j6�ԣkN>+�l�ϭ��]	I��9�x���V�=�%ZZ[&��ͱ�M�^�@�� C�6J�뫁�����@W^}�O�--���?5U�OK)A���_�@�4&O��)y��*�~v�[>�8_�m�,�)��b.ڦA����z֦26�@��9Svc8+���)?����/+}2~B��=�+jA�Z	��i�D��a{� kIα���x��*�����MЯ¹��g*���ᗴ�Jj��?�-�$H
�!$zT�c�v�C��ZMɌ�Ν��0���gI�V����v�_�$nxmp�_�3CO
�y���1�,��y�ŹB	=��A���f�5��'!���F*W��J�����~�� ��;'��%f�w�}��d���&!�z���� ��4DP�P��0gU{�8�x������~�L4W�j�#��qj�w�.ԃZ���:_���m��%�Q��ّ����?TH񂉘�s�]��Q�P/�`�8�%�ٕ���3�sʌa�����vG��
 �`��=NKc�u?G�Ud:B�G�%����t�0��)����
�v�XH��_%�e+�	F$���B}�B}L9��̥�p�>��&���q�"�+x;�,!9��w6��M|��r���)�� V����O��D�M�����P�O�-�^�q�ZХryK�b{�Ay0F��N.�3�}��ظ��us�v/mץ�c ��)�q�y�5V���� ����-�ަ6@���h�i3<�k�/��_�@�x۾�23j�k\%h*�E������4�#v�ף�Sq����U�t��
-���:��=�8���\8F��}"Jq.�o����)��A��q�m��.U��0m�Z����C	v���	4W�U�*���<���*�N~��c˚�j�ήhjߊeEi�N�W����[h��e��C(��~��YR���`��J�*���ewi�\�Z/�9v(;��A����G ��Zh��u�07�`��u�A���Xw߬87��OCsɧ���v�j�(���A'���W�slJl
�:ѥ	!6�ab+�F����(�8S��ad�T�O��s�ϙݝ�zS����A���J���]���w�TA*�	�QR��q��l�]>��N�KO�l�)�߆����j���Kʨ�r�%�����`��H����p/��3�V��wg[�jI�̌��������=������K��~aV���q����󩢋ȟbW3��d���߃���6���/a��+2�;5	�;�����1��Br��@�Ú^�4�ܳ�&�X��)�G���r�yW����E7�,>� �����f��%u깗�ү%�{16;_�5P�}I!��w�UG��x긴'���v~�D�?k�Ď�U­��Ǣ�\~�k��4k˅�!nG�ܡІ�:��2�_h���nL��N=5�<�P��b^�?���~_q���v�߅�̖հ }�$ ��X��h5b�Vѽ�"�a=���5����{��·En�BT��%/�C�c�v<�%����ξ�;x���H�j�*U��_��`�|���\cVO	It�'_���fE�9Uh��:TK:����D0�c�̐�E�.�#�-� ��T�n��%�l >Dhw��.���B٢�gBb�o��$����3-����Q���rd%�q�:I�,��R-1�*�
 ����א�p�JJ�����
�-*"��3���[V�"���hּ
A��r�>���{#�^�6��<��<A�>%���	���#^y}����#��?>q�vA��8�H!��n�fa���"�s��_�{v��5I{	ŵQ-���k]��b��H6}֨�^5��JD'��=�.U@�Ց��?v���Q���&���=�7����$b�#�勝��Q���Tn�D8(�ʊ��m�U�3r�Q+i,L��_/�r�Ar����zZ9�u{��lw7Jab`2	^�+��n,�jM����vw�.��n�>"�2H��46�VBڣ���0buE���l�s��P��n#U��hL���B�ܗ��ߞ�_��(��-������?冢b�USP �n$�ƾ����_ڠ���Z�c%]C���yFQY_��{�~VԹ��;�];���cOMt���5	�ݷ\ť�k�SB�J%�A�9�Qh�k�+����Bwɺt����\nӖT����^��v,q���m���N7�����E�Kؽq"���v��L��J�8��l
��q�͌�P��i©�n��J֠�H/ ���sƊ�Q~DU��6��q?)=ra{J��F�����CؐB�4B\��"�T�ө��m���mc��K�.���6��&x���W??��&�X=�xf�Ŵ������o\_=��&?���UuO��t��K��C�u�laȡ�9�qc���~�(�P����_����{��SN�t��3��2�,A3���/e"�I�w(��Fϼ������r��s��v������bA[-�To��=֡�&�����6�]��ҩU�S=�M_�I+@*���{�_��A�D�^�"Q:~0d�JF��`�X�M$})��2�i����j�B�d��� k����m�Vʠ���r�2�;�(�'A*'�(>'�N�^;v�2Z��X�qh ��	�0�jtw2�1�\��D%�}|J��gY�TQ?>G#vB����	��VZ#|�9��g���j�_K��k�5T�rbN��}����3�K��������Y1�(!f���T� Ў(���c�����τ;��u]q�M򼉾��~��{N�#֧�H!�H��3H�MAVd�C �����0krZ��N�&�@`{�O��C��Y�8� �o�T�.y����7��I?q��''�y9]�i�"%��o�Wr]�S����[ُ|+$��|�)��$!�L{g;�;�U͸rO�ك��o	�v�}�[-P��A�t�%e�@�R �E��e�+l�30��=&F)ց��\.��=���ZT��}�0G�6 ��%NN���F�g�4N�L� PS)�ѫ���jm��K��ܗ��O5��&�-]� ��i��]N=�z[��5G�@q���EV��F�|B�#�2~��=]|2P5��!�(�]�*0�R�h�
�ee�7Ւ9�:�q�5J�q�뢇�mGݵЋ>u��$`��c���Y�P0�4�`z&g���<���c���a�.qI��@J��x���
~��)?a �n� V��������d	LȘ�Ł�)�zs4�=�%ݺ��l[6��5/���Q�3�Xm���u�z�:����B���Ό}%h�ҥ�c��j�I��,��Im�e�If�\46�$���y����1!����-<^��m� ��:�8���[+�M=�74�lC��LK��tJ���S╟�v�oq�Q�r��l�M���!"Z�~�PZ�ǈ��JfR�|o�6�~�����LgQ�������͌w�VI��h��S��u3DSD�h._;�Q��T�K�@�Q��$Bb I�^��"�U��k��Q�>�/Z�(�m�������q(`�S?���`Z�hJ�bTo�nU�]�M5�>�n�%$��P�/�?�����H1��<�a`iy���i�Q]	�����VO�Sa6K��t;�<V�a����o|%��Yi���P�#����5uKZ�Lp�ܷ|D�/�����?ׇ+Wj+��&\kA⚲8礱�X� ߤ��^�~8����9M���K��,},�R��'��蹙T�$`��S��q�g>]l��x�.�Փuκ\�ڥ-?�b&��岓�I?�XZ�v���;�1�i4v �D����_�;�*�Y2�>�)�'�ͣ��3M�!� ��^x�:{ׇ�s�2�S�渽E�
���k׆���W?�5�|D�6��E<4jU�i�P�ȎV��"Y̡���.<���O����𫛈]3hi,��2���u����1��+9^,כ_�O��by )�_�+k�|I��,	4��݃z{�#�[	!���O��)����	�l�gl2F�ʬ��w��" ��t��_����]�+���K����'�xᯌ���^AD�g�M�l)K^χA�#���U$#�x�d�XK�ν�Dr�9Z�4��59ھVY�G��B;['sy'�ܯ���n�!������t��i"Uс�Ld���nOR^-�Bf�d0�M��Ʊl��@D96�T������)����f'៻x�*BѲCh����ʭ:"��@b�7��x��F��s��ڑ� Stǐhp5�Xo�L��.`�Vt:F�:b�˴e����7(ę1#���T���#�d���Z��B�1���s����ms5hp1�`nm~����Y`�Ƒ�����Psr��S��� ��q��"���C��ÖK\�7&u �U,jT0��Wm�TY������:���R����k�B�׾`g{�e@F�?虀���r�S���vͯj��
����<�{����xȶ�"��V䖼U��cN��� ��3;�ޜ�aS��ʎK��{����;��������1�>u��?&|��B�\,�ld+`�K��g�,O+'��$�������j��~��Y<�&��Q�tB�!�6���Bȷ.��$Z}����asS�ɡ/4�J�{�8�72�G���`B��p�:�w��!�����V�
�?�j7�6��|~�
,S���V��\3�n��y7��[����?�m�?���U���E�wV�;�T7�w�)`);�Q1D�r�G�]�Gב�z����na[K[n�w�F������/�Nr���;3��� |fw�W�uEE&��N��X�#�lg!Ņ�)I;�r�j+v-j��U]2)��2�y@���@���'�=<��P�U�X�&�b����xG���t�ha�k��o1�~���Q��fj1�^VPTxqt��J���W�����,�a�L�!����Npv?N�y�Y�Pc�J���b�������p��СGK	Vf+<�Hr�]��w�k�K3lN�	�K']���s�H��L0Aǌ*�2o�LRي�*@ ���Q�H[�r�`>�52hk����\E�9�,?���G0�4K���/=FKC��LHxi����Z.;�V8]D6XS��M�����_:u��̟w�/-�~�"��+���Z�Z_�� |�p�����)�whO[o�S9��Q�R��^����8��cw�p,�f�*]� ���;2��Hjb�3@ʓ��vAl(���lo��ğ�?��X+�l��̶.�|:C�Eo�3�@5�.j�k�K丁$6����?�	@��c������m/@F���1�����*a5g+ndw��ϧ�#�8>�7U�HZ�+�޹�?�2�a�^���SS����/�	a��Zo�8e����"ARk7.LBMe
b�'����hv�S�mu��BW��>j����my������^H��I�#�׼�yv<�wr��R�gn��%˺�$*^��OE7�O�2�I��8��nF�\���'{�!��o�����t���+�k��;@1��UQC�k��_tkq��~\QZK����^;&���w���N�Ej���2���� ��_��
�^�Evc�R_��i#���b{��	U���8�Z�!Ia�7�^�mڅ9-	��ULj�Ư�1�|1[�J\�򴰚3������!�f�����|�_U����3��O��NzGg&䧷��xx%�@�F=O��{��?�W�n��E�7V>t�k�?�lY�U>���kcA��(N�,_>�'�r�*#^c9d(&���A��=�1��[3hE�(f����'Pn�@�(Y�)�|I�`أ��A6��b+v ��z������#5�ӵ [.�gHp`H�Bc�AW��ޞF�kP9ϯo����"<���	"X~��<|�E�|J"*�L��NB���NQH� �^K|0��)֤;o�B�z 镩5���-Qw�8~���H,���z��Q,�SA`N!"%�!XyO����F޾���l�ɥg����^8�Ҕ2i�D*����gq҄鱗)
W��x��a�����!�c�'����^"BJ���ri:*}2Ew_k�uxN� Rco���czv�Y�'\��~|���\t߭G���L.�69խ�B<.H������NW���hc=��ڍaol�Z��A��߽�Ǵ������Ξ��;�6;D���[U�B�\fWf�g?h�)+G%v�c�u���6 MP�rt���LӤ����8<*#Q� ��{�ܰIY"rC�A��#��%M ���k� ë<z�ȇ���iw_.�̑}�<�_��4�iIwe���/�)����H��?�XcM�2p�f��.��U�Q �q����C<�38��~
H�36-�ˍjsq�aM0��������ã���RMƛL��+2d)jm�#�f�Pl[8��s�A!a~PQ���AZc��>�%�$0�v ���a
��!@ެ^�j.RU��|�6%<P������~7�],
��wwF�jy�:K~X˽!N~M�hy��Z>B��<2 (��!>H�ٹ��6�Pa]��Nj=����V����;I�Z/s�:�(�)y=#�Os�k��܈���=BZЧ.6���1ܦ��۩���R��}����%]~$b���Fݜ[�V��,���ZGW�?`���D$����Ys/i���lOw̓�X�l�a�cMg�q5�h9�ݕiґ��ܓ�8#ȑ�娽w�K��hn8�����Z's?Uu��s1Ѭ'V� �p>)1Xt��U�c��o!"' 
�J�o�xHWۈ�G�G�C�2>=�N�1eh]B�
볙�B�a�? uf�=Ǯ2P��+���E��k(U�]$�O�O��ך�чS�}���Lh�����忞�н���!���ڌ"sy[�X˓>~�9��Gʠ��ʌl�~�'k����J�؅=pG��A��n�����㖿��E|�"���5�A.v���V�^;�ql��ߣ��6L�s�C�d⩩]C��HImؕo7�荄��c���/e�b5U�27��Yk�- gX�QV��P^��h#�xޯ<��?��I��)zנ��WR�������D�,��s���v������+��
�Ò_� ��u�ΫS-�Dۇ��^�H�z�o�4 �qw2�,�i����[N|�7�<8��ߤ�9�����KT�S���'�(�X�9�s��]��:=�g|���tdY��k����4�Ӆ�&DKw��S�S��`;��tns{n��!1��`��ý��4�T,�T�t������"�^���$��#]K����_O�aV��i�텣��smi��ZR�2�e�z���x�3X�
��l�V��0S �ߏ���5`���s7K�C�|�̓y9e���٥�C��%+N(X�|�{�5��Xg�%��Ϣ#��>�����k�ݨ�N�+���AƣP�h�5������f�QE
8�TD�КE�}k��Dw�h+%�mį��+B��[㕞� ��F���ҿ�_h	�)�Sc�8��`bS���7Z3	����Dv���S�������d�Hj����!����\�-��1ƻb>YNXR}\��~=}?GZ���n�_�B���""��q�	���>-ðJ�I�@�5A�Nu?S�2��a��S2�d<8-�d��\+eN|I忮tRF{�30�9�X����i��3���#t��A.���8�� }�1�#}8ӳ����M2GQh�n��T"G�;.��d�I/`��:k��^�	���ߠ��w)^u Z�Ĥq�G��3�FJ�� �-�����Ng��&_�)>��Eˣ8���ߣL�Q��u ������w��V�*q7%H�,��e�Z��(�-�^o?��Gr#G��i��p������^���K�Ձ�T'|�N��8F˃ۈ�XH7�hĀ��t�t����*���I3U'I�Ӈ�-I���TN�m~�U��y��M��jJH\��9�5��X	�5�h���0Ǻ˞Z��J�gb\MtD�L`\Ǚո�ӹU��(-l�oƹծ���o�x ̐g�+�[8��X����EYϮ�`��!�u2À.�2�����Qv�� k�lG��ꍙ>�n"��ۭ���~�^%�8P�^��M]'v-v��g��ʑOEDr5T��v��%r~tY��d�H�� eD�2ʘ�q�l+8�oۑ.Ӽ�k�mP+��u��$��>�X���;����T_&��|a'O�v0��ŸD��PYt��\Ԇ#��}s�'A��$K����BX�5%l[�y�3�'��EԂ�kk�s�����ĥ�|�?r���o�Rq�`���f�k�m��m}���$����׿��9����������u�]�g��?I�v�*��v#�� �<�k�HU:\�|鎖�y��z[һy�pr�%��s��S���հ|�~��ik��:�8uG�n�J!<��⊍R���|e�ɤpL�b�7��\]hx��U�.2��ᛠ#2m��=�o��ߌ�>�^�� �f�t��<Օ�*�G�jj_IY�����~����I6��[FD��1�Ӯ���AL��7Sj��s�~<��g���cU�c>�#yO{�N�����`$	L�͓07����v����LN�B�^т��֙R �Y�x�wN�<|׏Y�F��h����=��W/]˫���3�>��B�Up�Ho|c���
梠v�
�����g9��}p@�DeZY��hw4��F1� ���.�_��	҄Gi�;ou��l1����us�g����&0TB��j��#/ld0ޠ$����tP����ĸmG��Ǒ^�Xꍜi���6�+W@����z:��W�O��q�8�h��X����R�-$��܀�X��i4#3���f��)���D��J|�k.�4���.A4�s�;������oѬ�Gǻ�L��<���a,�R�����6�l��9I�:����Y��8����֥�.a���&s�J�HNy���eD�`,��c��:�<ty��y�K�B�;�L�I�w4���Q�?���v��}����*���y�\8#z���w.G+�����=B�y�"��|QL�|s ���'ѷ b:�H����[�=�%��y&w��Y�W����^�i�j�`Cv*���tH�S����A�nI2��Ͻa�f���S̎e�>���FG�3��|�B�0>d�M���X�W-?�D���i0Y�e*���� 5�Я��H.�1h3E{��"�+�6��Ѡ�� k�������KjBIg���9T�I�v�0iK����Ѽ�E�h ��j�����Y��HU�4B���ً�t/�&$h��>q���W��^�2����=��l��l�t��d�-��4�����1�A#�ț<]�4��)���{�c�i؏)�L��&�-ҡ�4Ѣ�����0��c�
�UJ<�#悂��;B���
͎�\+7͕9��$~��G���C4��~�/�iy�V7Gc5I��J�BQ�m�����z$�.�GK��!�K�p�M2�_G���2�/Nƃ�m� �jT�0a&��\�^��Q�l:G��γ�¥i�NH�V���g0]	Z:p-�e+bf���})f਼��^es�U�]��鏰y�������o�S��4tc��L1]fN�Z�.�k�-���k��`�驻Mm��4����땲�`;~�1ÿ�m�Զ�R����3�z�C��:��ZR|�"��V緱�I6�) q
��Zjq��^)��O�w"(��}���)ʉ]/��	�f�@o�p�="��w����/5.���W@d�U2���=��q]��o�C^�l_�T�$b���F�ʡ�����.%��J����m����b"�1~B'���TFdHH�(���R{<p�[x�ӂ$���5 亍��Qn��/Ԛ�4��,�0�h�t�5?�H���f��wo��b����"�L�e0r�@���L�תm����h���?\����eg�� �@��nȈU�Zו����Z��Lۑ��@�,"G�;̵Hw]:ʀl,3,��-��dKROv����O1�أa�~�6�4��թy�U�1r���,w��:�4�4]^���p|`$�������ي#⩍�ė��%d�1v$�k���w���4r(��Lf�s�c���,TP�b�(�|�ߖ�m7H캈�O&p0�mI���R��eda��ۭG�A� R$J�x��_0A�3�D�`$��utdy��J'���@t+?�A��St���.Wp���E	��;��7�;��,��"@�s|���t�TMV�]�M����)6�/�l����rn�7'��J�N~,�@{��SV�ڎ�7~|f@|#9����O��-lo8�1Bk�㏤ٞ2-=��hB��:��p"�A������x⋧OOѯM$���EyK��� )
�=]�m
/���b��tf"�|�9��B��}�rKvb���O	ݗ�I���M���ӡ�h�h�r&�P<�?�6���8s<Q�rJ�Vڑ.\�@��>x��M��7�����m�C�4�9��¯(\�a�SVX�'D�n���G�Ls�xNG(����������*��O�r���������I>�-�D��$������2_o{ ��z�g��:�6KY��YrcDh&r��V�-��!S�OM�Te�����ŋ3+a7����ā[��Pe��b���[Ξ����Z�<[�]���(/���z7���8ɶR�h����9Ю��o~��!�i�k+ MP<�f��i�K⹮�z��np��=��&�WP6�͘�����<�j^��QT�޼���e��v.��܏BB6�{%4�պӥ�:�k`7;T�E���̕������ObԚw��5��I��
�O�����H��]��9�7]b�=��1���L9e����Nc�����}�G%�N�������{����<Ԧ	�\�u8��ݜ�jTԋ���!m�:1F��w�q@�L ����Ũ�-3sE��3&��H���|���[1"�B'n��<���cL��ݣ�©����sH˧)�}����DU��� �fH�d���徴T����Ő����7����KzX�4}�x���LZY���yx�|'<��@�d�~h���e�A�?�>���k�aϢ�g��[[.��㜃ܱ�b<~�1=*�&�;��'�Ν���s[/��v�����p9�	j��.L���\�s�mU���-�Ƞ���#R�Ҵ��")��X3��BE�l�t�n����a����{�����.1[:\�s�����]��,X�D�����a�޵7�R�E�b��Y���qՍ����w5d�:�9�e��`��\����9藪��@�D9ӧ驇kྭ� ٜ�)?�u���)����_|-'68y� ��"D�*V�0�,���r�������FP\[
q+��g&Fv6{�������</�ȟh��h(�+�cS��ŖW�G��*�=�͵��&��$��h���o,�uƯ�����7��i��H�w������.ܘ$7��m	��/�9I�sg��/������-^f��������ǎ�m��V��ny�\���������v��}M�a�ɶ�!9��7߮X��/2,'U:���A��,�g����ƝAjj1u���3R'
 �{�>��`�ѫ'�=Y��g����e�Cz���i� ^%�rz�e����ٴ}�/�f�����C�x�i�ݱ��9���WxE�$�/������P�a��P�̥��ٚ�u2�܌8FA�����ݕ��	gk� !��^�Ӌ���Ќm�U�ͫr���V���S�fQ�>�{Eܘ�����{�����&

��� z(L�T�)]�kCb�39-�ަ�`}��$���=v�
���[Upg�ܢ�_>��PB�ķ�&am^�}���]��@��o�R�/�2�KS��i���k�<�c�%�fTX?�Y �M�ߙ���B?���l�9=��K�����`�d7���0�6!�Fi*����_g)Y&�0��9�8����׻_�+�-��X�u��F7�*�����6!ڶ�Xm2���n��,t�M��\�,E��r�-=��ֶ��pvG@Q��e����!��>��C�T�3��J �h��C����&P@|������ƥ��f,�U� ~��_�����d����^�1��_�d�֏l��E��H���M��#�����z��dF�9[&����Ev�0���1�5����|�,2�F3���c_�D$F��3\Ⱥ�m��D�� ���n� ��\�J(�!9d�J����u�X�JQ��E��&$[!�Ώ��n���Py r喝έ����Ά��A���NPo;�obt�+	Z�⾫���c1*��g���9 ��,����m��L��uTT��`���шk=�!:��y�wt�x���L��yLYZ�uٓBE�V�I��΍S'j�3��qKw����Y��}�}�����h��*MW<��rcr.箊�����[�v�}�=�OP��(S6��3I^9�""��Q�%�g'z�f�=>���>p��s�d0�������(�uA
99�~�Xj�T��>�����i����ߎ���[,�<�Af��Rq���$.��
'��F���� ��7�٩�lJf���G��7���Fj5��?��nJMGU�7�-�i���A� �ӡ�����q�N4�8�!��O&6�@d1}��#��-�	�p�������G�* �	W{J\�Ѐ����-�~\A��4t��2��:tjَfD��$��m}6�t��f�H�]d,W��/�R�`��W���Ph���/�����,aH[�2�������1QWl<��b�����h)z|4�9�+5�T��$ߜ��\L�3����,�P���[./�q��=��|� gҩ���	�՘X/G�����,���F}TAB�=��<�%Pΐ{L�����%��q�œ8Fc9�n��cyh
U��_SV#��T.���2�%i$7;"��}3䫔"�G�3�����'n��>��3�I��Oʾ�f��Ad%t*�X��zf���d��e�w�3�ޫt��"��()%���=�|C���,>'������>u�� ��X@ٵ����S�ja���s�W�g��qL4�!K�!�յ9�cڱ�\k#Z ����$Y9�o����Zw�[Ȕ�*�x�i�_�.8~��-�D��,�<[<|y3���_ߗ��F��u+mzEm�2�T
�k��&~�2�"� 3����D�榲�KT���GC����0�*�Y�d�\���Xp� ̀@^�)��A5}�Yl��ӦK��(�e�Z�������7���̀�Gx~(]�P�B5�V��:.�@W&؝�m�L^����9�>Oh7�dwy�$��.�.+�>P]��Hx� ����-+Vgj�z��V�Xė��s����Mf@��#F�2s�k43W\��B��o�8��_�<�9P�u�b�x��C��.!^�d	m4�o�G0����n�k���5"'��Ҭ!|���o��I˪�ȅ�vTB�!xe�/?���3���%[3��X%�8�O�Aڑ)O	�3K�ޕV1���
��J`OY ����B�\9���z�=����w�kX߮��Y�{2��Gi�[�������]/h������'�gLPp��|.\�}dcO��㡘�ڠ	uݏ�'xI��dZ�'��ȣ ��TH��o[@'�M�Ow��97�\L�^��-jI� ��PsΌ�����S��Z��ސ����e�@ԍ_�X:ȯ��t ���)k�~�Ԛ��dO�k�@�A+�
%����e�g!$jVCF4ܲ�8�ٝ��{��"�Ɏ�����<�V��}J�h�l��.lDP���]*�\A����#��e�:c�xq4,��+��Ed��� ��O�}8wG� �2P����C!�}n�Ʌ��qX�9\EHF��tP�5�f����Z������� �0�)�dm�^���N�;s�h#H_�x�0���3 ��l���<���!�����-�D/�0�Y�i�+�6&+R���e�O^��w�H����fk�W�7�'�I����� �9��
�����/���@Y:�6��8��z��X�0��4!�ld�^'��&tv���U��VV<��N�+n<�T��HGo�/�<�`��mi`�b��Ew��_�PO?��r��m�W}N���	C��r��pl
&s�H*c��`��;&���!� g���Nj*_v�\y��l�t9w�������MB�	��*E��[���	T��p3ZQ�¶��d<�k���Ϫ�ᑇn$��j��|w=����ِlbw�`4�Dߡ�/Z���G�����_�n�ùO�,I��(��i>�!�(}Ru=C��)��-��l���H�G����i���W���fX�sa_TP�y� ˵�����
�#<jm8��A�����NY�+	�Ō��}�W:<(���;��T֝ez7?�%`��G���쬃m�Ҫj�F~[�ѝu�0��D6�������_���`�5785��I����Ҥ"�Nۉ�Fϸ�+Zy�!�+ƀwQ�ێ��"�wK�Ĩ�\ö���z�������#�Q���8PL#��;u.  ���I�کJAs�U�L�u�K�P��}�%��ޯ�cTu�­b����T�{d}�ıV����'�y��.0V��>�HZ���S���b�&�#��X`f�f����H3��K@Q6%4�������i�(�6���*�.(&�C��P{ ���Q����2����*�"���9���r��kD(�=���F.����m��=�_q�w%����XT4H�7ዸu\Rv���^wl4j5�0��u�t��w؞�%b1r�!n�[��\�P:�we�����[�ݷ�F��F( g[IIs����~���c[%x�_O��	�ރ�J��k֪�@P������kx�����ߞ<�x$N���%�?؟��!k����A�^��]ETڍ�.���k�����a��2g���W�sT�f?g�Or7Q#K�pU��2�
qa�1{u��s�'��%���e�)�~!�ke"��ꎷ-��N���GB	i�W*�L���~���1�P���0��c���|�4M���3��F���6|���P��.��3O8�v��	�4����[���)��?!8�V���3@FR��x^#!9��ҽ@������C��]�nK�&�A����������}���_S�B��N�����_#�ً���z�G�Q;m�`�����F���7)5NUM"�8.dΣU@/%-���]5�p)��#��$v^2aî>q'��P�	F�ݥ�O�K�H���'P��Ძ��N�?��\��-�����Sx�"��_C�8[���������f -6�jo����nй#�,������
�e�Z�D�y�Ȣ@_`3X��k{,ȍsы�q�YN+Qob� ם�lUI��A@�\9D�K.��n*Y)�V-B+֗��g��o�˶GD[��(a�B��f�a�8tnR(gL�B�z�?�g8��K�&�<��om�r�%Aݺ�v���I��P�r��	��C���ޟ�;#�]��&�X��hԷ�
p��1M��J�W8W��0=��(�3 r��0��>ڐk�)�D�.��U��.���K�9ܜ1gF0��6���h�2� p����zl_��2�E�;��ie��R�@~Ǩ��U���������~A�d]Z�g����Ul��kuC/�'���<�X0'<P�č~\�}6���
�r�%"��llZ|��ێ�׻��p�2~����-/�����*^~�ݶ�Q:��r�E���oX�7������ݟBv��~n)n#�§=e5��~�P�b�vt����[��ڒ������-	2\B�4`�&���
2@�5S?�ʙ�\��h��a8~�8p'����w���;��
��@ɶ�A���%�$�����T\��@q�̞�.���D9����|�q���2�]	�R�������2����7�s5YL�.X;`q�,#Y��M'�
��3+za�GLzԐQ�Axqs,!̃؀�fti,���v�.Su�f �˵�G�uqh6[�c��Y:3`h�6M��ʮ�[�ZAzW�[5X[����ii��w�������O5�tI`�����O�iސRĀ����ʹ�}(���C�703�	I�Ei/W�X�n��4���Sc�"��Q�z�d8g�	aBu��6(��粅L��	_��I0!ƈ���c�:EF�tmI{sq�Ń
s@�)YF��[m�q���I
�G��2rY����@+��z�����؂����j7
���Tt�y�`�fH��=��EF��0ۧ�	F]�8�N��ܡ_�A_�^�U/la�h1.0BPS,X���Bu��̂lpa��Sl��vr��sH��X�NjA�K�9 Fo�ۇ��1@ۋ�&A��)�T�p���Qe�'�ڐ`\/��Xj��M���_1;��"p��#�Z o��	��e��.e�:󏱨��fk��M��
��F���ڟq/Wiڼ�l�4#�W֝�q�#?��J�3����D����j#���V�w���bB
>����Nʫg���AP����X�5'!l[�bM��5狶,��R�?R� �M������1QCW	9����
XF`p-L��@��͸��r��KR��i����'�e�`o�!҆�4��v���x4�I>�DuA��P����j㦑YsW�\��pK*JhƎY���$Cf�g�jA�0w�M�)�%Bf�R�8��=�_�u��w�v瀹t�l���QS���"+�$��l��=�i��Z�A4u&��?O��i@������;"i����#��v��EL�<�l�E[�r��"�t�@�Ͱ��V���]�sc�}�2�q�ӺdsH��cv�3�3��D�s����c�*]��Y�X3��nir�1�۟z��L�$[��TK�\k\��D�g�br����� �����aS�.��UmWtX�
ԛ�v�U��9�Ev
����~�L|E��֙���+ �v�5�^H�\L�9�N)�(AZNu7�.�{A�9`��B����7��#괆����[=���^���u��t��L־��|;Sk1�^A*��b��L��W��̎�op����8��J9�҈�?{���Ai���+���`zc�c����Н#:=��T�8��w�U�B�I��*m�3~u	�e;���Fy�2��yv��zk���[�� ��]]lL���_�NI��FI��5]u�=;D�<(�(��[�3=����y�������ESm�B��a�!v�b�۱�|J���l '������%^;�3!�{T�cxl;����'!\�4ov�S �2
0S�s�u���E��/�꒍a�ٝ"���(��A@���c3L��X�[s�	����I;W N�
��6*��<���={�L{(�w�]_��I�c�N���k��j'�Ǟ��7�7�t�Q`�WB^��q�Me�C��ZCj钛�·
7�8�w��"���x���<�<��pے��W�|n��_]�J�8:�7S�Ѻ���3d�5b�3���"w�:K;���/8�c�����g�
Q��S���0�vpޟ�1򔭻��f�V�5x�X�����J.'M2�ᷔ�p7�G��,@+([�f�d�A�(t=�ܓM�W_.�m�)2\(M,���������Z�[�s��^L�n g��.���1�����Qz�2 �Mۮ|����E�*�n>�SR�h�K��sPM�I�m�d���e`��4t[2<�D���cC��8_��:!�זf����F�Dn�Pt�&���� *#Na��P�0�0��l�����\��c�v���ظu���Oꆆ9P.<m�hc�<`�P�0d71�&�s�)�@$Vl�	���8�'ٛZ��+�S�zw'���s������G�K����`��u�*�6d����ݛUZn��{�)bc|V�D�bQ�$��G#D�.R�S���*��F�T���x�ZDA��QʛYص��b'#C0�+&�?:����@�n��z�Gw(����e1!d/�7&^�@'��3G���l7׋��^YM�s"վ��OJ�w��n:��0�)�:��$�d�W����H�T��O�Z@����gm�v}�hi���a�k0�eh���'ӌӯJ೦oE !�Ђ�pe��aCn2S"y5�Lǔ+&Y+�j��&c�IzO��?I:d���P*��fVWqR���!+�M�K�sN�<��]+�7�o~�`oa�o��� KU�B���a�;�qs1Y �#��~I���²��h!��o ��*�2|g
�(i�{Y����J};�w3
ߣ�	P آ^r]�i򜢁n��t�f��HV�\S�����k��GBŔ���:H�l2p�n+$�(�h,8ձ>���
����8ߜ�%���x�P�FZ���M��z\�Z�\�a�#�x#G�L�8B�X)9�t&s]�4�i�T�P}V��߲9�%�Ζ�!�=Gp�8)o�vɅQөt�q�P_��?�g�"�&4�u0�U"�\�]�L�/�ӳ��[g�ZD4���ό��<1��:$:x^+�z��>Ԟß�M�w��9�/�ϸ����V���P�������,�¡�8]){�V�������¬����8?��e��̈
	f*�E��<��Qq�n���(ʱ�j�L��X��Y�{�PǸ��� �.���*ʤ�Ս
�8S�G�������s�^6C�T�BS��g�A*s,��5��%��K������=�3Q����D�K�く`��2����>؛�'���K+}��^�uc�IR�̧!���X0E�������}��p���J?����IKo�DLo\�-XR��*��&��B��H�*������MH��c�y��	�Z �/c,@2�{��IO�R;<|���6_3��:;�6�J�`[*ϩ�>/ݻ�s�i�4�;��lV�_�N���k�c�a�'-=H��U
g��\��� +�����v���}����w��R�����	�OǬ�P�Z("��+�#Y +6��TR�2}�e�ʭ#��Xw却	SGóh�����p���&LW�����HCF�����+3P(Y@e$�*�� �]֜D����`��=���[�c�np�P�hqh�bY��yw�;@9!�k�m�x����U��)n�ܽ�f�����u�d2��=W�|f�Vb��� `ȟ��Q�4�ʭ���b� ����st��g��"��5��Z�B����r���Ь��9��؂��`-�[�'4��.� \��~C������>��
~�o��(�U�$�K�<�A��(��X� �C-N3yb�\�����	�&�������:�@���s�_
��rE���i�$� ��]��n�[}2�j唅i�s�v76��~�.�je�.4P��y�#&9P��lm����4�Z%{: ��hV^r�4�j$�p�n*i�F�hj3��]�

�?��,��?���)��1�g=�cJr�}s�y<�a�<Ӧ55ޓ3w�a_��9�	��A"vp�A�_4���{X �6���Xg�M
�ۨ`�:\�eQ�&��N�[��I�Q>J<�I��g��<��u����҅��~�`R��M���<sx�x��#PYl�W�ǻC����UՒY���Kp;`Y��@��$3J���ɵ�� ���;:����^��)jKe�*ߌ-'�)b?k=�V\&��f~~NC�m�*s�椔��;�q�%��?H7_��x����ER�wӠS��bf�xl��z��
�R 1���`EG�i���RO۱Qism8`�gA �Q�������2x�O:*N��/���4�k�Ϡu�w#���ZhnP���A���]��pF���p �W�S:��`plIq��8�W��t�b�?��V�g����2�L��4�{�=3;&�;��6L��-P��L/%�7W9�V~̅�����1"'���r��e�-~t��i�0z��IkC QrC�rC��^{��>���T	m���u���/�>�R���qY���8�A���� =�'}߈!���K�I�`���Q$|�Q��)�.��sS�%�v;j`gu���?��g`�����I�莈/�%�\QAXȢ�M5�J �����������O��׺Ø�\S�9 !k�D1p����S�Bf�5�3N�@�4YI���� @T'��H�NH�1���Ip����{Mr<u����g��k��#��NѭUeu�$�Q�m C��LeC�*K���i���<���*\�ߗ�:޲J�}��� ��s�#��&�,T[�6yV�✟=��h��ѵ����t�X U8�NP��m(6T���Z����I�Ԛ`���~jleft�2�A2�%��	��a}_�cb�xf�
d*YB����-�3=��hդ.57�/��^��݇��+r'��T`�R=ͭ>��A�]��:a�{��CC�NXw��_���HQ�!Ә��z%�� Q�X�{i����&9��ˇ�j�Z{��ʗ2�N�S�㔗����oD2J���8/kBL�h\MK�*�|��\� �P��R��0r#֜�-�6,��8�;v�lb0H�-^{���\ئ���M�I�����Sn�|�n	"��HL)G�&]�I���9$�n_Y��X`�j�=m�-'ɱ;�}Gt�����hp��*X܁�H���a�Ə)$��02k�kЙ:4q��N�x&�⤏o��l���A5v{�����}�M�G��F��������y�2hV����X�7��;@4-���s�+��z����$�9u��+L�B�yK,"
���#�g߯�H�#���MI='N/g��x��/k=o!��\;����0~(h�W��X��[��`�O6�\d���q,����pgN�R���a���羴�-�,Mo���
���J{�����?�D��+�0�Ƣ6���d=˶\�hBœ�Ӻ�i\�㽳�(�Y�����a����T.��@,BE؞�3�0cjK	�#�����4��8QJ#;ȟ:�J�.��E��%n#K��C�c��Q6��`cG�;)�
�o��R���J.N� 4C�~F�-�(9O\��>Y����R�ot]��+���M�l��yn�z��C����y�{Q���]E�XS1\������ GlN��j`���2�-�ۛ�$9��O5⹲������`Fg%
/��9����ݳ�:55��E��N�bߓ�/EA�����>�緻�\�-_X`�A��%���*���)\d�t*�]Or}����*C6�icI��:^�z���r>������`��wO���Nn)��,.*���͍_�!Uej�94�	�	�<L!��.����O�˦�R��p�A]��e|���̛����m�+P�9}���r�i�^v5^Q��&�����R��f 6��W��,�	:>��Ջ�lbic�j�1���(�!�}��ʡ�561s.�ʲq���{2h��Խ��.m۶�z���#܎j�RH�������,�@r)�Q���w'��B�lp ��?��h�҆A�@n ���aW%7��k��Y��u�MH �V���Q���2a�,b��$,�3Zw��G�8V.,V������ɾ�5`K�ю�B�\���	�U����6O���U���^�ue(�nE���r�{
�J˳�	��MQ�yy�[�.n!$�f� �T1I"��;Qm�J�RuY~#���b�i�+��s�P�m�}���w���Ӻ�<:Z�$�<m� F��v^�ַI�������U��w?���cȧ����L�d��_��FO���ҧ��.���T���۵z�l({���X��~� �B��SQ�� �����#<�-��B^zm�H�;g���N�:m��J�P+BT��L�qɪک�9�[������l�Μ�]q0P��V9c#�^�-��T�Q@��H�	ou*�L1ap3{3�۬x�vHӺ��;uZa��+���ǀ�IAڸ���p\ ���sm�ж���W$�ucMv�[�`�����l�TB����!�߭�_�IY4��x��,�ŗ�t��:�/�k�K+6q�y\E��NP�N��go��:թf�Ĺ��� d��ҽ�x?�G�7R~Ü-+N�-�耩R��E`i��k2��[�Πҏ!��Pn2�;̆�&��az��}�j�t����;Ǭ��~L��O{���DH!g×��Z�h��<�y��`�2���]�;�;j�y�i�kPr�$H[��p忈�ꋷ���F�i���l�O�R�4#U��`��12A���9���Ր�?����#tI�^l�)S=d��#���L��KG��К�*�_B��TP�	����Ȱ[������0�(S��\E]��Y"o�$FA����X�ڢ�/箙>G�	�,q{Z}@Ϳ��O�=!}��Z�Z�)6�g��;���'p�N��uZ����Ĺ���o;�'ܤ��vܢ�tR�R��q�*}��
�AquM�j\��ڡ5/��ǉ��,�Z�*�#��h ������\�W>���څ=i�AGn�ə1��O����	^�b�L	0}���M��2�X����fD3֛�Ȓ��c�ԣB��:���+p$��'}�;�X:2S[����&Pj���/�;>fҽcv��W�\�t�F2uTkW�`LU�YM:����;p��&(RƄ�4�ڨ?Kro-g=g�l�����pk럹q%�m��r��6�'�����9X��O	|��&r�]����rÑ��Q��{,nۥ�x�6{;�y)>㤤���eL4-�ϴ�����@����ϼ�{��E��#�R2�:'�N�>2�|�,�G����#j�(J�n�0|���wxv�)����L�+�xQ����HE����v�(c#>tԳYg��-Z�
!T���D��ßܖ6�����yY֘�z�:����9�<ѽ�HC���9���OIC���k�HA�.gh��*O2�w��X�d�r�� 6ۼgv%�O��37��T�����[���Pwt��=R�_�^ª�m���Y��%�k^�gu��U�htu%�Z�UGZ�IkD>G��@����d�q���fE��|82˦�+\vd�7g����y;4�ϯZN�@�H�ng�.�pӘ���[���[�B}��jd�`��J�U�6���:Mj��<#a���i��B?�E	Խ���0hg+_���P���c�_ډ�,�Aϭ^gz`���L�ڼF���`+�]�����w�ؿElmv.�H:������$�9x�I <FT�������N��2h�����kk����v��"���T�f��FP������cV����m1�M�#don���)�o��A��*��~�^�zQ��I^�������0�0M�K��F�h��8r�$� )��&V�jՌ��NH�м�I�`JI|`O�AQ,ܶE��4�m}��&N���G�F�b^B���)��]��$�{*^�1��-�׎���� ���L͖�i8�����F�d�<�382�D��G��ο�m��:2���o;��3M�Gƾ5�ej���1��z'���C{���!a�̡�)���R����dc��B4vb���|�F��7+�s�#F��m��YO�~eFgC��>�;$@�=��T�(0�67d!�h]��H�P�N�L���g��9� ��Rǒ��
CP�4V}-�Po�%b�fY�#�Lew�%�Eoͫ�YJ�ח]�%Ά%6OH� �"�P��@dQ���E{�$=X�S�BeP��G�u�N��<�������s��
�i��$"�]�[N����?&��%j��T�k�cxG���+���\�oh�a�,��k�����"�#)d��6��lG�%:�MVX�[�|�^#���7]�+��ߢB^������[��7-�ț��	�F�=�l(�P�P�4�D��r*��a�B�L�zW�jw�#+����p���˯9_���z/ ���ٚ|ڪO�M|���`�$2�$�	èea}�a��ۗ�c�vUU98y��+��r�G�+ٵ�mf�iM�'�.���Kw	� ����5(����P���]A�e%�)�f���P�?��KŶYFyQ��>��e*G�)'��E�~�DB�=Pn7A�gԖ���s���`$0:�d��q�J���nߎo�.~��@�![��J'�̿��n�8T$��7n���� �tn����b�n!���jG�م�Fh���h�2�|���DX�����W�Z)��^�k7ثٿXǼ�/d]�n��=:�{�^K#��C��g��Q�e��|{��v{��\7c����ۨ�u��U�5j�ҭ�y*U���|�o?����ZԤ�
z��O�����b��|�8����X��a+QeG�P�����+�WM�����с�mc{�%̀r �s}��|�<4ͳ%�t�D�*�<�nH�b��l6[)�y9<,�е����ky�7S�d		���xڳ��΍&.Mjώ�\!�A#+�Y��ZBa ��V<��Q�f������!$FR�J�rf%�3��O��0�j���j�����	_��Y��a Ԇ�^i��] ��$�Y�E����BO�K-;v��5��̵�\.�z�䀅�� �E���f�e�'Ģ�cUs��O��DM�J�9연��$9ܕ��f�u��O�J�h����4���>��:�4�<�J�'�n(J��1���={��RW^�����{�;j�B���果)��7�PU��A��&�����\"�ۑR����[U~�P��+�ng���"�JBS��tL�v��Ւ�P��K�����{L��6�Dn��$������/l(KZ����J�^�9����f?�!Q��":��+5�#N�~�p!▐�z+\V]��W��]w�+��H����4(u3_�=��S�����C�u%��կ^�B���e�F�}�0mh;9/Z��	d�vk��+	v�W11��C��U���0C����4~��,nS�(�
�/O���}�Q�>���:`-�����X����������{�ku磦t��	ƚ����@e��*t�Mㄿ8�Y#�⩼o� B�dU�-��	���=�h]~��:��k�h!#�W4Ey�Q�`�OBN�$I#�Z##�g�Ӳ�NE�q`��Ww��N���>-���u�w�N����SYk:0m�dJ� 3���l�Z�pKRh0�/��.�n�2�+�n���k�e@�cr6�c:e��R��I��=���_�r����U��^�;�( /� ����g��;��v�M�|9�)�8��[ސ+&�"�U��;1'p�D�@�jSf'3F4\�܉=�k@Lj=����sV��8�e��#�:����jsS]F ��ޫX4/�C��5]�/�p�i�1��c��_��+���DNO�Q�˸L%�P�c�9�y+ia`�~_�꼍���pYԸٙ �'A�'¥f�=��P:����Ǹ%�1�d��DC�`ڵKG����ZR�-mz
ҕJ�J�#��lI+MW���g}b�3��%�xA���ᎋJi�"dr�ԩk/t����`q�L�𢖛�8��"���k�!~��Bh!��VN���a]�rL��U�4=��R>8��)��~�Ѫ����Z9<���@��o�qʏ��3�;\LL�������������:i���q �@�~v�;F�a>�f8E��i&�}��#�ā��`& "�^a�Zz��
�{�^�|KEhk�t�V� �?�Ŕ!�b���p3'
���Y�kniis<��,�`���v3����1��ý,�TH��o�`�-�\I#�ky���Bc�|F�"&y��N[��+3��}AV��-��*���|R޸�drr��E&$�,�̉���2X?h��#���U���B2U��7��	�Y�!ַ%��\��"�C�%�^��Xec�T��:����9��9����JT2�g���b3�t�!w9�S��d1erqR0@�4�\�<�&ݙo��U�>�Og��*1��ezc��g�ϛ�]�a~h����dZ��$ʯ�9�wae~=_6Q.�ǌ�v� 7S���7�ܳ�-N:�%/������ �S�'���Ե�4��OL�B��Ta����ܜE2�&Lx!��� C��F�֢(O�>�Г=T�τ�~X?���+A�Ðtt�V�),,�>�jDJ���5L?���i�I�:���rC�x��}!N�RR�?��2h]���-!ؒwS"\A�'z�o�Lv*i��8adXB�� L� 6��q�!?�)P9�l9�m�-Pn0ҕ�Ç��cb���[�0L!�������V��C� ��u��z�ʈ��RT6#�9� P���eK����&d\�"��Uc���*��,��$*��1�4/ڟ���E�hOMJ>qX�QWh�\ν`�ؚ�ڥ�9���ۮ�0�+��́��FT�c/Yy�:zh�3����=2��q:£,i�&�"n�U�҇l�ܚ�lZU���XÃv���>�P[e|^�:�ؖ��uC"'�"I�&���]��J�2ѱ��8���y���<�I��l��n�M;Q�Yw��H�ܚq8<��N#����ް#cb:�: EvGK� -��I��a*�����J(��� fkd�W���lb�zA1Po$P�	�*1.����1�
8��l�ʫ*Vg+0��9긂�7�N'e{*_�o��\�ѱR7���UJ�[_�������\�����N��d<�U/�@*�;>IKq�-nc��r.̃CQ���m�@T��J�gQb�Y�7�u��sZ��R,n�|�FtaO���m,��R�뛠�g �x����*a��r��F��SUKh��>?�~��Ԩ ��x�a�S��widz�y]�9۵��K��f���m�K��xgW~kr`=JiG����# ⬀����D�E�0�q}�]�z�,��)0n����P�3#$��$������ ��+�-J=s�:��Bc 4�.`�BQ����YB��c�����Ο�0��y�	��H�Z����U�?V~3\�u�^�4��Y�WC��m��U��Ƒ�5��vI`3P.v�mS�S���,�(��o�������N��ƵۆڇN�w���(���u��^�dk� �I�x��R�
�^#?�؍�����?�q)���u�V	��p�zqx��x+m�/�S��uu�
�����l?e�	�L�Q���C&K��s��u�"������ŁWz��V�Nv�A���R�nF�V7P �����
���z[��U"*��Tkd���%FE�Ɨ�7�'?���	=pu�}�h�}ZX�£����$�Yn ����倚�����Ѱ��N_��IE/USN9��:}�J��M�:S��}�gݾ���	'�^T��2}�Pk�๚�W$��.�����ѣً �a�Oc���W#�"��w�T!v�?]P��j���&V\5�ۂ��8=���~9�N�[�����у�{�&D�t|�f�`*�#����9V�4Hk�'�s���֧�){-���%OΚ�b��m�Q�Wc�gܱ���Y-xN�d�1�;T��ݗm5K���y=`*��J.a��de�b�F<IխS����Q���|��S�E�P�P��q#-M�ý�l����{`=E/[؆DB�U�3����~�R� z�Oe� ی�����\q��J�3T��q�j���SeH(YV��J���b$Mw��vn�B��e�u��>���הvu��,A���k�%`�^��"��h��QU#Btq�϶��< ����LlލY����0_�fE��?ŗ����A�^{<��ۊ�4�cT�{l��?ƥ��v��Sw �q�z
'0b*T���C���� �V�^�X	�IS�Ij�?�_��kڿY����y���}�H�^V��ro!"�x7lpZ�꟒��hh���ۑQ�
�q�.�k��-!-��.e^=�ۥU�88�)��h���A�j��2$�{U�tzJ]�Zi�^����x`�)f,���N��)�h$�
��1E���AKPz��!,{��h�|��*���Mf~տ��6�?_�C�w��i �Nʜ[���w�2��C�$?!p���V�� � ��v�6����V��"&���;Pkd0%�
 ~��x�8��䗣��l���eg>Pk�m�"B�o��O�gw�C<M������Y��{6S *{Qk8�R'�҃�,h�(����|�{���a����q� ��d@V�E�U4���w��q����ƾa�0��{��cx��:���hom�oF�&��-/3�w1c:�]Y��N��zm�ش�y��KSd'fd��\WFL�WI�z+-%����>,�r�N���Z�$�Ak5��@�\�S��b�W!X���:��25�g"��~)/)��c3�a��$mq#(�Ȓ�	,@��z���܃-�KAE�u@ �M� �,:���51��;��W��3����}����-O:�Q�jA�.R'�?�72�n�_:&����G���������`��~��Tۮ���Vb��o-�����$�Y��=��nTS^Qf` ͆Z��Y�J���� ��Џ��AM�Ex��Q�~�1F���C��(��zФZ!��蛕��Wbq]�҂���(1�Oq�	˄Q��$���)�\s�;�tO2�a������x���I~��6w��;.�%U"�K����2&���.���¿_nX8�I�`����P����������z$�C�r�4g�lå�^edN��]�M� z����2�\(����?"�8l�����>������p�y�\T�A�l�t5��P�s��h��tNϒ�]v�
��Q5?�_5.�GpI�}��G��kӒ�����U���s/ԋ�M+���a�-�hk1�'�V�T��c�N^�#��B���ȋ�A$�%,92o��1ӡ�x6RF��L�X(1��]�d��C_z���<إ{�sbC��J=�`���'�K�d~�xm;������a9$��Љ��$6p��@��fsNm�%�M0����^�vk`�г?�)F�������^��e@b�{ҢZ�3����:�H�rǫDK�՗DZ��o�er4-!'d�����xDND;��=�� K�k]m4��EI�p��ͅ-��}d}��UW��Ζ�Ǹ���x{�\xuC��)b�|����O���[���̯��Npo=��w�㿁��ިn| 2= 7=�t�/�-rl�);{N}�z��ŚM+��I�D�H�@z��>)���4V���_/�Ϸ�~�S©X���(��b� ���
N�n���\�EZ��P��2�mS1�v�����oqazm}fs@�!H;~�wp��m?�z��0r�۬+lsa��.OW��pԁ�}L$�8O*p,���)ʦ������f��? 1�壥���3;au)'�0�Βn�M�j���y��P�ZA��v�ڳ�C>��F(�D���^Em���Y���Bi0`P7e�^�����2΍�5�w
�$+���W�������%
����a���-1��Z��<59�����3���E���}[��mȞ���*O�fIdj�G���7�8ŉY��4
H&;Ɣ�+c�rؑt��z� T�ĵS��ѓ�%6�|�%�Eq{���V����D8&W^5Q�j��*�O�?���[W�
�m�i�U|
�_�Pv� �����j���8{�H��l��D�1;�v^�g�@����?l��9x�i��'��H��9��f�ԛ\��#rеZf&�_yA�lGH��M쳌���=D�܏�a8�=Rg$!i8�8�E�F'Y��G��#Z�Z'�x��B��DP���u���kT�"���	2r�<0sш�:�&�%�U$��v ��%�!�nAd�"��hM1�{�;<�A��4���/~���nK����F�k@VW��6�@�t-��lT[J	�m�Q
�j�ѯ2�kZ���������&"_�)��C�����k�ex�32�C�iL��Ø5���s5�W����fs	��@~�$�*���yh�
���-E��x�#�4���q^���m�p�P �������EA�q�𶀓Uȋ�Գd4>�eXw��Y�2$x8\tC~���y<�5E�L9ze��OBCPA�uH��.\�ƒU/H�lla	�p�9�:h�|�� ��� ė�k�+P���ni Έ��[�`��_D�{@��?�LeM���?AXX���x�7��?�����f�Nj;�E;u�3U�L�g����]�f�%�������ٕ��1wMZ��v��7���(m�ss����S���Ҧ~��qqVQa����cv�"��̲��t 9�=z�F��.��k,��Iv�8���4va�X�`���L�`G�>�v�S�4��~x�UƓ��ݟ��bE+M��*�h�J�O�v����Z��A�6���������^������?b�@�d��AN��M�vݒ��M>t9�
U�r1�y������d��)y޳��sǄ˜c�g��%�IM@RR�;c��ʱ��J!�E�� �w���>N� �HGJ�^*P:��U }t��b/:^	��h-�ӣH�Ɛ���g8Wrp��us;�&-J�}
��`�L��m-��U����~���Eq���ǿ���Hrx�M�l� *:��^�ȩ�#��xTo�`�a)��_���S[rD8��j�o`����b�/u�VfG_j̎��|U3Y]�͛U�1mdTVi� i�5G��V����$�m��"V7%a�����%/\���c���.2>��hFS	}Y~y��=3�?����~��]상W�Cl[�[ ��DCԣ��m�3���_�6A�M>�#:�ox �8��\qq��Ō�dߞn
>O���U✨�!�������k� &up�ѥ�q�����O`c82�V��Sʘ����JB�D�xJ��������ƺ�]K�{$�ł�X�p�����B4?\.��γ�_����3���z�h�f�����7Z���s&� . 4�U0�6��YpGE�(�i	M����J�_��6�('D�q���ͫϥ%�/�W�:�+]��$�y�@JH�`/G:��RJXd�� ;� V1<rͭثp�&�ʖ�>w��+��� e��U�!�6���xq�f�O� �k2^��d����~���?:�Rg��͖6Z��h5��2|@����;/e�EY ]�v�B�⅏-�7]��<?�t����=�R2�S ��򳶎�ڣAc��r��M�{�[���{���߬�X���A�kih�)���a���dN�' q����n#J&vjYd�)�Q���pwM��a[rw��g0�"=�h�ب�1�}YW��]n�.�'�J?�2Gέ��i���n�g�Ƀ�P�7�K~y�6�o���P���xUy$�!4׃��ba�\�^�!���ק�g'����3뷿{�_�Ot�~N
�I���3��3@ ���!_�����U�i�lu�|)���L��y/�o.��k��u���IU�e�F�F	$�N���$-��N���O>G����}��ƕ��f�[*$nb�6�^R�e�K~�:�'�C8��.��Ǘ���ٵ�y9�,��*p�1����C�ZZ�3Ap�b��@=?��ɬ�_<�����#'nqZ`҇�O�������{�5�;���_�+gJF��l�Fv��XioD�)2��X(_ �$�.HX4���CJ��B�~�b��1
��CtK<�	,�M��K.�t�dW��{)��ND6��hzh1%T�w -�%�p�P&��٦CD ������m������o�߳YY�/ܴ�Br���ՇB�m�Is�Q;�[��za1X,,yE��0�T��2_��u�-�l��Eja�7�=�W�eL~�0ހ#Heԣ�!���$l!���\:Ε�F����1𽚌k��,��,��;I�
+[�4L]�t�y]���$�?�n�u����C�i�9���Q}Jk���a6�dճr�)�h�[���Ne�$��>:��;����l#qI�P�U0t	b�<��i-�7�\]�6������L�{մ�ؐ�$'q�͜�N��@,+�=%�v�G!�����;�sD���b��A"�xב����c���������Bﻪ4������;E{�j$.J}.�/�AJ�2�9E	"G�bo�����Ө6hf$�����Vd��GS����ؔ�X
���!CT�����K�e�8��>�����Eb�9�߿�i��)-o|�Ę �]������H��d�ޥ��4��A ���i�����?���	�/��RB���R��
�qO-1�M�a�>��z�3�_����xA����̜�d�lO5ȹ��_�t��L������I�I�����%�Y�,�X�#�\U�lu��%���/�����A�����aW��X*�hq����;�C���|߭Q ��2V�L?�����4G�ᰭ��%Q�S�W�k+оӊh���^y ����D$6��?6���u�W"v�ץ�����L����1��\��z����_N�I'��H�K0$6�*����չ��'A�4d��H����&�����:�����K�dW���8� �AD���oG{�@����Y��A��?�3ۍ_��o5����f��HS��G}�6Ƣ���텇X?��$.ߴwN
�����d�S�c�;�ޜ�L{�ۋ~<�Ӛ��`G�Ōtm��@*�L�v�"+�9W������QX����Z�`G���l����;��n)�z�8J�W���3*O$ӿ45��y|�8�)M-S8��)��@��a ��sd�4�i_f��O>��V=����7�0og�_|QV�GU�*�}��1�����������p�"8�ܯ8���в��­S;���=J�L�ƾE�)��R25W���]�V�r{,�_A�|��ӊ h��\�O�n�H�.�g,�Vf��q����@���e�y����EM+"�H�Ұ�;e+�r��(�,Syz���U�n�L]<����b�ù@<�T���`��x�������]2ֽ�miq�/�j3����کD(M]V����w�4�]�[�>������JQs�;d����Pː�1+k���}ݰ�����L�K�D��IҩN�Rm�H�y 6{��MR��ʍ�WP�V#!����YC��I��엀jx�`;�2� �=0��uY�5��[Ea���4�8����r֏�%�n����MR�Z�'�(���sL��:DV{O�y��+��Ya��g�ϧ����8 *�ގ�TA����� �M����&B�sW���!N=����s��h4<{����Iut�B�X�(�ʏ�:k�*I��Q�L��љ��A�����.�/���	W�^����-|z&p6� ��d��c������u��A���0��$3$U���q��������%�����T�Z��׋1�9hZFi��E��g2S��;������yZY����Y��V�%����sοAj=g7<+c�R!��E�
L��9�t����ud�1'��$��Ռ����}�RUI�}�YX;</ujh�|��*K�!"ϰ��E�z�wje����p ��Eq��~��9�$ ��4n�ɵX���=��	�8a��%�r�4ʼ��eF�|��ab����`�a�	D��|G�����>v���ދ�ec��i���TJ`�r#����$�s���5�$� O�fQ��a�#[���Q��O>'��N�~6%�� X�R�6��q|�sÝ�Qr�[��Q��c�y몳S/;�����k��R�w	�
&-4��?ӽZC�o��"�u+�2P�C��a�f0�J��!�d#�!]�}N�Q�hD��:P͝���N~�+n��S�5�١jZ)�ֳfr��
A����#ĸ���Ay��fT&���aC����6\s����o�b�&��S_ba�ƣ^��ɘ1�?��x�'g(W��`-��%�;c�ڈR
�q �M��X�����֮Q��K�\�-�=Z���;5d�t�{�χ�n��m\�DH��"򎀓�!��}b���D�U�(/��A1�����ӫGr,sHG����U���F,{�-`�Ĕ�S�B�2]��)�wJ��:��Y���|0���19��m[��߈E�%�i��;񖹞��ʹ`��>��֣֟��9�?�<�ClH�]�$Y�92���%�O�����C����T� f)�v��lsôqm���	��ĖӪ��!p�����dP�x�	^�E.�v�,4V����4�	H�k�MB�nkR��$h�vy��1B��d��o�9uJȿȍX�N�rq*���:�F��(��y�W]e���8�>�$P�;X$=�vUX�Y���S���7�,:�67Н����f��Ic�^:��j��$�Fbc����V�e�	��Fl
��ʗjH�[�W��[�V)����@��'��|��H�`),�?�٧)̎4�4H:xۜ�Ջc����k�@�˰�JHV�%���7�l�d	^�J(�%��h���05�j��Х�a�#C��!*0�ac��L�uH�FЦ�3�zN̫:D�&/��lh�8���Cd��ƫ�����V:�yX<_�� Hʣ��.��iQ���M�F�A���;��E��U�(�U-UF�ϸdw�d�գ3��$�=w]�:��L�-������(U�љ6�.!Kи�}��nn���������(���[[�p������J��0@Q�f��4� Q&*Y9�"@a32�=F-�֠�F��!�L�J;F��=�y���·��x7��ý.y�|S�L��>�cZ{n����
l��AUuP��HN��aL�߆�T�ԃ]kܦ4N�HP=n����$ uѭu�xhK�:�p�=Ӗ������C;�	��m��g:o	L �h�)$3V/m�n������*D��Dܑ�~%r͇�S8�9��xt{���(N��(>q^_<�A�xA�gTT����?S+F^h��d����>�:�ng��� �.�&���?ڋ 1�] 3��\{n�4��؃���j�=�qc/���:�خ|��gQNMեqR��`hT"�z4�/�CZ=kQQ� TiP���yh� p���t'ɴ�*?n�$�Z�-7=#���6t�3�īb&gl��_h%�������)9l�eI�7w�y��y���#��lsS�/��<۔X�U=�:<�u� �ޭ��:�~o1;]j�����"d3���,�	��+�R3%o0�y�ë��k�>���S�ߢ��M��tӈ�u8�arN��ł��Dѷ�y}�jr���=:G��M>#~�]��j,2��6��/:4�Tw��2�D���TH��E���E6�{�P렿i��%ok�N�i,��Ř��<�9�M"	L����ĸ1�J:�(�bJU����>�`�AOљ1�4u-'�>�߻��K)(	'���ꛔZ(U���&쐇I�xG���t�y(��a��묃ڱ�m׃�r�U�O"v��q/+���s���[l��R/5P#H��g�XEE�X���[5����Ώ��܈y2��N��gl���ԇ��^b���z�E���uq�n�M�m�a-)w����:)$(���J!��,��.K�FK�Y��ү�v�ɛ��+ts��#������#H�x<��[]���I5nX@��/��듚A��荃����LE�7I��ș�A�����K��:�1�U�0k�dC���ʟ�X��A`�s�h�QY�C-|�$��aH;��")�iC�Vo4����r��1HU��+FE�t��-!tz�[�H�f��ad�}�@�u�}V]�&!5�?O+����*{1���+J������|��QF-���I�Y�G�؆bM+�W��N]xvh��O�p��J0r�)���]��=�*V/�!u����.�B[���k-䮯_.�����%E|��Bp�ʊ��!z`��O	�L�˼߮ԗ�+Y��������?���51��bkV�
�<�D"����;�K	_�m�S��iAx
������ڜ�\�E���9K}V�Ι?��u��z5���� ��id�y��1��)�5x�����]�QmBg�[�����/6I��	��8x�J�&`�fb����/�R�D_W�˅\5����C�Pȕ,�Q�9qc�l��^ֵ�g��:N[�n�W��X�u�%��2@�nD?̘3%G�$����{�,�� ,�|��}9�8���R�_�gh9U8#�cL2�M�_�<�L����J�1-B ��lV���ͨ�b< �&��]ݚ��$4�-'6���o�WO��KUYi�b-��wQ������)m^-X��k�86�4��m����LI��e�!j�v,"\L�D'��E+�o��~d���2�98��y�e$�6=�>�|l��h�^��X�m yC�NѝFy_�� z�񟏔u'�O�����I�"���<�)��!�l߉��x_��Cg���ϳ�)Qf��Tz�i1�4�����f��ߋ��Ґ7<2xk��󍡰e&B�!$n+si]��0�j�#�XScSM�^�"�V@/S�DI����i(�D
��h˫���H2C<S嬫k2T��%�M���2��!���X~-Yi���rͰ �N�Ȑ���{�vQE���(��:{�\V�۬o��~@�)/���^�}V��v,^���I��nغRN�S�ql�a�..�MM��7��v��Ǭ�����^�b@�3�o�'h�	 �m���'�]T�E S����:�S鏄��LD��-%�X��x5H�S���d��7��VN��/�ֵ1m=}��;�Q�z����]�0X����n^4�U����d}nE�t�g!��R�hƯPJ�s����Hpd)���x��:5k�$.��=>���z﫿��[;~K�!�H�<Y�PЛ ��;р]��"2; ���ل�i��c�c�p(Wc{�rjwX3�` ��p6��reg�]�x��T�(,]���;/y^�K���<�P���}��:�1݆W��(i��+��6~�E���p���D"ҋի�t��(DJ�"c�F]�cn��{ Ǜ>i|�S�<��5���{.0O����TZ�2����9�O��J��.�&�1��U-��S,6�ׁN�^�#���~v�o�h$=m4�C��Ek�}�
zHQ?t���W�x��j�z�5��sӐ�x�[2#��s����AG3ι�:���F�������t���@$qY���Χ%�����GvAf�EO;(�4o�H�i���Na�e��-�sд��}p�+�jЙQ�M�&T�%�0�ʷ��N 
�����,J�{�59t6PP�6�����$�s��>�!���j́�U���r����?�L^RW�=�0��{�S���"¤��o�w΃����~�!�E���q��C"-bC|�Meߌ�TV��n�zAc�Exf�A���D���OC���viU(���|���6Ui/HV��3�A|�u�h�/�G%F����`$�w��q2b�i�}�59Ĕ�gV�3�
�����R�V���R�u�ƆT��5]ۃ�qڋ_�Yg�Fw��ŋC)d��]����h���:+T��!�	9{�d�����Ȣ諄�d�%��<1�	~��I.�Y>�
M{vҔI�0����i�"�ߙdw���M��y��@F�t���st']��͝��@��^+,4_���RZ��g��D�)��\L<9�������:e��%����M�� �C���@��R����{l�:�ĕ�7��n����Qz}t��Ŭr�A$M�y����8�`��a���Cr�2�a�Q���n�ʒ��{?-<�[*��[r��_��ޔ�:3Uόi�f�'C�ʑ��@�{P�d���)ks&y	}��ʅB������C�@0��� � �U�#��CE�B����
"�h�^�A�Dײ�����3T������7�"�3"@Qc=h3�ѷ[�E�p���{����o�
�K;㮊�-wA�AH:&��������$$ʱ.������
�&S[���ʸ�� ��l���@l�3=�Ay��Υ�"W�(����<A��vֈ,}� F�f���RCo� =��\����S����In����xm�q�$:����=5�}����ч��＆�v����Ӣ��J�XՃ;@�j7�Ѿ�uI�����;~�}GR�V}�i��j�;a�*+Yޑ��GlR�r�UnG�ށߍ�Q5�Fn�t��55�!���,�ڵթ�S��=�d�#�5�W1�cA��2�\I� �XKW������4�p]��.�$�0�j���t�� ���>��I���9��N7EOK��To8���L�יZ�Ct`���+��x�ݰ_���hѽo ��*ƒ�޴Kڛ�5z%Լ!�iE��M��P;��vv	�B���?�$��{��b���v�Nt�Ap��I����_g�gfF�4�q��WfAmǧI�e����0�Mѫx	�I�r�+�CP��:ö|�h���k��C�\��]�r�Y���e���}`�t��'gn�\b�Mաg	h�f)�>�}Ah�������dn �����[��6�ZQ(Ć��M?���5ʏy������Ox�����k�pΟ���J����t�H�m�s�6���,t��,N� �`�L&��RX�3�a߾�7��������Nn����co�i�1��X}}�tWh��-tj0�n ��F���[��a{	B��z/����rc�O�� k��-�6�H[��l=��2��mg;�Q��m���j�4O���	�!�P�Jn���������,D���195>����=*VvRȭ���$�npJ{&BƜ���T��f>B}�P1�sT/Q ń�{R��\�L�\��ݖo��T�i�����04ŗm��-+��!�S���?�Fe�I(�[t���JAͶRjԂ��n��HZs�r�~��C��k�|�Q���3 ��K(O;��0z;зrFe���.%�;&$�� �	�dʠ��E�ت�oj#�p����-�+e-wQU�(�$�&����	1T��p:� 5-8y8W�qrк
��(I.����3H���]�w.�H������\Ъi�.�j?5��=⚐#:�S�PR�d�@ۆ,]<z����$�}�ƒ��O�i�%�ח@��OU���r%�#Ep��=m���V�m�de�&�B����`I�D�R9�ˮ������HNRħ�^�� �4q��T0ܵ�s|�g�s��������z���ǵ>2�@��E�I�-��f�U�A0��
�����/���Z�eB�ܐ<���}�9��v�fu�V��t���qN؄;�@�.�V��k�4�⾵���[�{(G`�k��;�JV0rq�{}�t����V�W���s� 
:��e���c{��o�3Gg�n#k��̌�P�>�o��&���͵)��j.}.e���I=ٛ�k4/be�_@Ǉ�u<u�c{�k�� `k�r�,�RM.�V c7O�K��_�1{��u�(^U9F���Nw���5���ж�d��:@p]�����> �]���:|�uB�e|���7]��g��XZ�է
D1=����h�<�6ߴ�,�j��r�\1������X������P*��"I�>!�z*�'ߪX� ni���R�V��}�����"ftS��&�X�*�B�hbf�����E���$m�+����9�y"J��(%(4�Ñl�}��V-m� �V��W��)F.\{�!:�3'���|u��ڸ�n�2��Q%�F5�V&��Tɱ	�0�`��b3���,���ߌ�	ę�@V��"g��6�btҘ�(��5όu�A�֪�	#�-�(ik?��)Q9�*��M-48T�� ��N%gZ� u'�}�Y�bG�uy����"���!i��<�vgi"u��I�+r�/����i�n����33C.�I�n���ʰ��8$7� �����Us���I��g��4��?X��V��.Є$�笁�P_IC��ҎQ���y�}w,���'�ˤ��P謍����Qr�C�T���(h%�gX����A 		�ѴnFM�Ŕp�;h�{Z	�5dOW�g��s���l'����?d�Q��<�t�V�z��=��o<$�^zDI��G��dlz�sz���;O_�3,��(��]2��!CN�o�!}��k6�,�)`d�=1��:Գ�G@�n�� ֦��xx�.��#��nX`�˧�
� Z����bq�g�@��Vd˯�?�p�Y�?w����I�ڍ�\��%�1�u��9H�a�M������G�Y���4�~�b������ c����|E��EQ�s�L��	���]�����/9_���S��A��$ן2�#/_"e�p6�?s�5	M��"m}&�o$���(@v qZ/���� �\ez%̾�Џ@�v�W�-A��+BC6h���s����^���M�d��}�P�ꖭ�7|
%�J��:YGҾ�u$�Vo������T�,�˪�[��$�f#�WB!K���<ǀ��,�dw��q	UA\T��&F��ʳ+�$ޘ�6�+�&�0'�I#�X*�`̱ �c�*�8k����*�L��J��a,6�	O)?������n��Aƺ�[��п8�]7�z���9����@3]�k<���}��1�0�6�-p���Jg+1V����D/�P9��N<�0R��,���(L&WJ{z}Bo���m��^@���DIbaڈ��3��|� 	yVc�W14�K�4`��6�P�-u�,-�q���?򋣑���qQ.�vzkG�ʩ@�3�P������^�><����j��@���]����/�;3p�����1Pt,��)��RB�2څ��E�\��#����?F���\�Q���J~19��%ћë�o�@<�\^�p�>�n�$K�m���N���P��O�s����b�`��'��I���)����
:�\c�5���X�B��=6�12�5{���PS�Z�!Yff@<���6=3I�`'�����$���_li��ɳw<�\��"Q�����U�������]��9�%���2L��i��In윏�J�YqIq`ֆ�h��q�++X�<vyTB�G���J9�V��9m��Bz.�X��l#���B?�,���G�d��W���m�|�`Ы/nv�-���a	�88�7h4�L�V.Qڊ����~Ar'Xd$�HW���sM�h�6P�F�9%��Fd���$�w$���*�e����@���qQ�Ӂν�^>���Ԫ��=��nv��+���T,f�Y!X~�b
0l�@L_�2�Q¯7��ʑ�=^!�K���|���ر����5GE����<96'a��)�	`� �J�N�cP�X$��w�@:�A�L|ɉf��]�#$�J��{��_$�9��L�2E2�t'u���L���vGA�����	����Z#7��vk��PZֿ��c��WnaI�a�6�Z~K:��C������⸐�1�`��� (��aq�uտe~i���j�/��\���¤R-�|<	K��<�;�6u����~OШ>UZ��T�l��<��~�L���3q�KWI��ö�@%S-��������3���ב�X>^���������q�^�U�0��\��m�A�.�4qK��]ez�z����	�ܲtֵ�曑� `�h�J-�j4$W[qE���m�Tb3�i"�g~���5�t)ܒ�����G����>J*& 4V�=�U#";�� {J�DtZ��?-*1Wȶ��x8&;\@=k-�H��`}���ѳ��XGGm�ĂyJQu��y��tZ̈́�;�H�Y6��{�e�-ˁ��鰥 �I+�^Y@�!�T�*@SB|�5f�i��Y�����vQF��w� C�Z9W�@J�y�Ya�Z^���硻��}rN��Y�=
���a�^���Am��#��Б�!�	k���c��#ށy������,H�L�[��:��Ȳ^`�?ke�":t~�Aߗdy�~U�rLǲ?�S�1��~�3wh��AU��-h�%�����mS>��=.b%О<b�O�X�T��5��E���j�{8UH�R��r���ߩݎ8�?u���8�����b�W����f`l6�1l(ײ�����.A�m8ݙr��U��5��8���Ő��(����]$r���0K� �ř�X���Mw ;�Yܴ�yIo����ݐqƃu�R����o��Fy:�(���\l��^��X`��Y2)�fǛ��02����f�[�y��� ]���+��*�-�(�mQ��ɑ� �7�D�B�R{�>h��x�O����ݔ����͉zX9G<"���]���跅]�0�(7l�$�(�:��\�)�Q��J��7�zc#+��u�\�#,�1-%u���p�೎��^��'�P���	���R1��d��4���8���jx���}諶
��˛Q[}8�<�Ƭ��"�M���)�;�(η�U�Z�� w&C���
�1�yЧd�|����u�@O�Fk� ��|���h���������99N�:/�C�;�t֍��34���蘆��v��u�E��Ujz���1f+CA7�H�W�A"�[쏇o�3(���]4������T��Ԇ�Mrd�$Ѵ��!��Y��m��P�����D�/�s�<dp���Ȣ>�=3��n�_��:���M ��!���S�"*yO��� ��U�|)��uׇ��@�u+�ɑ�w���)�!չu��#E���� W�UB��9e�H^)��֎-d]px�_�*]��F�^��W��!k�����p�/�ޠ'� d��s."MA�'���J�
��_z����FL��Qϣ��Ň`#`�����'o��ol����=�`e�-�����:l˹��,4	�����Z���3�-�EO˱��O�n5��%�aQ��f�aZj��e�p<0w�q��IK�Z?�(� ���ͮ )->1��bğ;����̮�ͽ"���䕭��P�5�ŎK��/���Kb���\���j�!}T�:���f�Q��)�P��Q�r]�s�NLw����S���N��-dì���1�{6������Mi�;D�CO�>=�����ƅ�d�E����-�#�0+jD�ެ���=~~�}�����.���d6��	lOO���evju��x��,+o�a��{QK���9�W���`��VR<O��|�g��>�	�s�]�/���tO5��(��D��=�8&�pT�p7��kP�yf$*�JH������]~��-�o� ��3�L��x�o��A�Vd�}�B�efn�=��}�^){5��g�'<^pPCI��"SZ��SD�q!9�&�Mb�s��&�s���A?�iy���?��&���P��PC!z�{o=i� ��]�+|2����֋���zR��j���S�V����/����08���@mx�y�눨U�8Bg��p�L/�FZ`S�V�,N._�H�n4E�ڠ��0�t	}<B4���ak�}��F~I� ƙdn�/6��؆��E��":��ƈ�(����^�hڛe�e��Ф׹�8��t9��y`a������ [Np�#p�O�K3���y�r!��g4�cQ�ĕ ׏����҂��}���%����T'��/�OJW.tp��	�;��U6��_�a�Z��F����H������}Tq&�����?�\��Dg����G�-KC]w��d�e;S����7(�-պ��Pؠ`_`޷ 9w4��@�+bsq�3מt��7�.�����L�.���fD���(?w����j�U2#%��`��#��qj�i��qr P�[�x�MѰ2�jG6��o����kо�,1��x��s6��.�P.D�ޡ���� N˲8oub�YA�R_v`�X�D�g�%����OEhdw1m���ʮ��oB�Z�q��*ݝągK�4oW�U��[���V����ט��{8�(/F.�����pid	3<��]b��-T���#\<���8��3���	g÷�|G0�3Gb���E�,���-�]���"�XH;XG�gSJ��C��E�/bs�v��W�����
8hp�b3����f�ɼ��90�[�hP��s��[����4/K9DÑ}�m#��D^/Ͻ��Ԍ�0�=��vϦ����k���qR$i�:f;��Y�1j*���N(�B�7>%�_����Ό/�9ҥ�o�rr��o��un ~���qe�{�ěA*�>���'fV�@g���͘�� &H��7-�Ȯ�ɡ�)�ؘ�,k�����[ �5m�9}�{��r�l74u̓�y��s�;�>�);�*��aŝ�p�r2�fI���r:��\;��F]�ui8�@�܃֯�!UV"�`�A���%w{�܁!Նxn�j�4�M��� CG��j#f�()LM���+uf�l�����4{�"�Ƿ�u>���ע�y
��d��*"|�����j�G��F�(��z??,� ��wG/i�7��û,uҏw���Թ%!��z[��Q�Bh�\�K�Χ"V����`��Kˡ ��a2�9F����i�Y��C�~�)mv�n��?���2�vPFWft�]�"'����]L�c��FH�O�]] ]!~�<�))2Ro[r��
s�[ݑ#�K�o�O�U�<�Y�z���
��\v����YZC�j�=	��<����L���O��C���ANp�߿�hx3�L)��
Y��p�]5�H��5�48�K¯�;���hG=�V����o���vy�L���Jh�U.�b�|c��g����%J�!q�"���b~����)Ĺ�F��Tൌ����Y�㈓DVEbT�j菍Pq����V�0��k�o�X�X�+
=9�Y5�MU��JǰV�O"���hїNP�V:�w��z2�zQ��S$0 ʓ >�1r�4?@��%퐬D�A9?�&]�F0M�t�1��^y�?h�m��e1|�AvA����l~�������O$�.pd��(�������l8�&���8�(e��-�D]+7���	�2�t�DxX���l���n��s[��g�˖IҚ�Q�{�uN�%�Z)�ϐ�SN�k��eYv?X< �[�U9�Ci�2�u��=}����Ɏ�P�i���f}�5,i�Z�<N/I8��0�f%�$��
��-����ۄ�z���ŗS��b�2�aQeө����� Z�
ٻhy��T���ۣ3�+���οi�#���fǆj�5�l��'f�	g���7��AE}Y1�T�(_��	7=��OԏY��L�(�s-/���Ŋ4�����!�ܸ�i�a��R�4����%]-< l L�'_�
�0]MYJ�(,隂�������Ѡ��Ď�(��|�=�S�W+���v~�����E^���f�[�˅��T5b_��*B����*;�d�b�]�c�=y�"�u�B�����O�Tl��:���ۭ�I�Kn��2GN��ntE�Y��t�D��&�23hr%c�{���᧺��%ӥ�Bֆ��jU���i�7���i{��G���@��dQL���ܰ��^�Ŝ�P��,�>�6��NW�5��iq+y���B��,w޸Y&�C�`O%SJ�5��e��I/�Np7r�p�%�H�1����PTo� ���.�kA�Q[	�g�&�(��3k,�̘Gb'܅d+
�~\�s+�N
�ā*�Ŭ�&X�06�ɼ�)w��(%�e���i���CR�yJ��' ޢm=��{�������O���z|��#~E3����Ά\��4�t��/G����p�8����ޑ�0�� ���$t��',����p ����M�l)O��g0�����IL��w��\.lk��`|��Ղx@���(�w�\j�oW��ƶX�$z��W����iE;����K�7u	6�	K�b�C<f�Q3��>�.�ؓC��V�V��o!"ѯ3c�g֙XŞ~Ւc�C3ܠMG�@�o;s��4.U$���p�t%����ܖ�Z����X��V�%%�����M��xv'�{��|-s"�0�?)���BΥd[�r1.����=��rթ�\T�u��_K�/�a�O�����O-u6=�d���E��U��9�˲��،
d�M��� ���#l� �+��a6�ES|��/�`*~U�X�C'g�j�!��*�Ɨ��zphnGK%䃞a�%���sC y�O�DJ�T�!��v�� v�־��Uz&[E�@�T��+*��fQ�a>A
�O� �w`�y���N3�)Oԇ�R�!���il�"!N8O�=:#X�|z���v�
��&����5�w��4�a�4���L_3���
h�nv�L���|�5h����f�6�f�+(i�nOTآ���?���B���V���p���Q��'V��j���V��-u��Z��ĵ����t���5D=�zW��S+�bopE⺼i`W����N�p%������.���t	�P;��mW���EհF���Tm�f0�XX�h6��k��0�^�cA�i�xe��H���$0<G��
z��ܧ��O��N]���~��7�{5:4���6���9���ڑ�l�Z��
��ѹ�Q	޸��D��2[��^>�6X�6�_c��8c܄�{G�M���h����\���-���a�{�c7N����a����f��F? }�lIީ��d�H̥� s��3�d�P-:-t �k�a��U姗�F	�c>ϑ�=�b�#���F�,?R�GZFm�5�V�Ȼ�1Cus�_{8��2o��vq��ۺֶ����<E�YL$��� 8VU&Le5D��� �P���Dx�D'�ȳ�.���FBlJ"�����.e�e< �Hp��ͳݟ�����ܛ�`�a_3tS5�>�|}��4)�F��˖�x*U�ٞZ��A�cm�ѡYJ
4�"z�Լ���g0�J^�]U�T�
�!�S�I�G���Zڗ�S���M�T�^ŚDӫ4*��;:��S۟�v�Ț�V��j� �>|��}/"{^:������=MfU!�C�R^����AYU[�c���"�PK�bK�V���?og4}t�t��d���jDϰ���A�&1U�i�A��yk����	CB�Ћ6��-|�p a�u����V&_���&��qq�6�↪V&Oz��3��Kܙ/+�P�7'�P����f���)���:�
4U�h ��k�0�)��r�i%�P-���{�����=tݠIv`�������~�;��{r4?��Ѵ�1txDX��S���(U�
��	 ��5�f��>��pƭ���썜FQW2ESѰ�A�f�S(S�Ǭ���nd�� �m,'1�����f3't e[%��cw$���{�q���ƹ~��~"r����);��+�b_H\�l��щ���!�1&�S2�9v+��n�|Z.wC�.�՘qΚ�n�m���R����z6;��b�s���`����o D���k.�\l�UǴ��[�Uz�W�4��Q����X�7���z����K d���v<��đ��I�"�p�wP�'DHi_�U²�KsُZ����!@��%�>eF�]�wB������J30\��5?�J�G�ӭ��.PSLy�0�P$d��l������FQj���R��$g��%@@��Y��LW�o�@���8e(FY�8jpj���mBq4���tg�������ls�
����4���L���K6&acw��5;!�{*�E_�Q� ,L�����A@Zx���?�6��+��Vݐ���ӆ�%���7E��D����qm�)Hq���i�r�Sk�vW�!o5����-(��V'��zT�h-��{�%Pi�T��n�� 4��f�0R���H�)��o�V8�_�ḯ��C����9~Q�p��ֿ���6�(��.<iH�����}nxc���O�qd�Mn����>��s��R��E�L$����"���H�$��ʬ��VG�@}�~r%<��9?�(~\����~H�U�K߄������"�Sy;�ldYD��Wp,�v�f�K.��֘E�"s�`��4y2���m]m�/E��ڪ��]�½Uլ��g�՚�)'�8��ͽX�P!W���(*:w��������V���F�̗������)bG.2��FIm'�o�tAZ=hk�:��D`u ,��V���K��������l۷�b����jv��D�$uAc���I:.�(PI��t��~g����0��`L���N��j).�$	�p���a���y�*9�c��|I�H���������tď�m{�
��D;sty@t��Y`�u�}N` �HZ"����.�ŵ@(: [t����4�aM��Qz��׶o%�<�cǦ��m����"�r� H��D��?���!\�)P"���׍a��V��}�H9���cRt�	~_�v�ȸ�a�1{�Z�)ޫ�M��ՠ��		��c.�aǂL1����$����1��N�p�C�F��D�)5���SP��ٰ3���m�]_#(�2��`' o����R-bu�.��-�T]�F�����
t��R�\{i��.�F�"`>R%���j5j
�ܑb�vb��{�ɵ4A/��9g�:Q}$�r5���͠�sɉ���=���:9�>�b��w��c�6r	�m{WudQĮ���w��$ ���=ǜ�W���aY���������zI9�g�K�p�yM�����.<��)���<�x�������I"Y���x�E���,�m�����(�Tr�を�U�]1_��3!���f�Q�=G�$������qp&��}��� K7�q��5 ¢������6�I�N�'��k{Hg2*5�����J蹥l-P��Y�П�58ҫ(�qXWQ�f��@֪��$�'�rc0�Ie!0�R(K�!�;TO	;���W����Ί�{7;��z����M^z)`�BH��
4=ZB�0�5l
<){��4���`�|R0~W��]| K>�
���V�V]ě��91@���#��/�^#�"fG]Ӓ�y��r�;o?��ב{y������K���ȯ�ͻ�E�P4�q��^�{B�X�sJBH�JH����m�a�+�+���C�C��wUՉ�^�n#���������X `P�BG�*4�D��LQz��>]��ং~���!^Ɂ�p��Z�o���9��Xq7Ix�a���	�-خ��|�!�"�	)����-�Z���[��� r5[�*K����|�>(��\M��E햗�i�J[�6�$�˩�%���JPL�
���hD�l�n:���5�+�V9�����V.�ZCŵ$yF��Z�T(I�9��o<rZÝ�ْ�U6�����U�vh~�L�*+݁b 9uG5�, �X���m&�j�.=S�%�1Ǹi�?(��{���(GT����H�����J>�b���KUM�X����"軝�(a�8�=��J_T�������)�1���	^��h#�盦+�8��BF�
$O��H]����\[#�qeO�h%_I��@rӄB��� ��1'���(�xTN)�5>�x��V�	s6�y��̇�+�@�d��&��"I�P����S������c{�}�M���C!�+&%]����QB�6�\&%�^�|�&�AC��΅��%�ŸƼb��6��pR)"Cs��g�4��A�r]̐:.�D<�i��m��I� 8�� 顈�
%�k:�<�f����2y�h3�61�g;��y#��kT��Y��䰒����t=h��G �hX�^���ɶ�jY�L\�D'��j�w>�1�s���Mʘ"�q;�z_����\���z���<(s5��T���k���w�����a�|^��1�5t��W_���[���_�p�>(��.���?��b�ҳ�W�І&�� x׬����ޔ]���\���}�>�]���!�Ґ/A�3��p����V��߅����)LEv#���� ��?I�X���:���z�DL���0�U�_�=	ār��T˄\z#������I�d�g��z�c} {�51�u�[ɭ�t�Y#����>W��-�G.4Om�Y�cj��w��\n�b/P����Ou�skɤx��� �Z
B#J�؂����F�����~�Q��à咡�*��a'rg;�����k���)'Rܪ:��ݭ] �(�O�.:������|/��
��2�Nƻg\Ѷ�mv��ۇ3��ВA�7ߏu������X{j>�ݓ�o��@���骛oY�۔5T�T���L���X^J(�Ϧd�-%^ Y��DH�9�����?�<_/�ǂ��	d\��Zݳc�s���]�H�B�5y��%����k����K'Rd��������)��~�n)*zkrx�0Y4=�5�!��W��]�]9�)'h�y�2P��v���[A���9��/�R�vaPDF�~�ᒚ~Fr��;�W�}�E���Ɂ�Y8��C�u�ƒh4Ȥ�o�p:�����mx)�s|��/9f�W5e��ـ־�1�Q!r�a5wҽ��.� ������O([���]V���Q���^�[R������C����H?w����&��4�աy�*���qXq�Ԁ����ͷ����C찉,�o�"v�#���6C�g�/ ?#�ۺ��D��d�U	��5.?P�Vv���x3���r}��#�ܭE�=8Xw�*sKx�xs�
���"z�q!�1up�2sh�@��d��Ĩ}�Ao��%�	W�2�5�uj7�*dg�׿���Hj��"@-ɕ�Ե�1��9�'v�T�m��A���+���aw�2���{F����IӞ^��,z\�|T3c+`�V�
\��gJ:�4%�=d�9��IT�1h���+��ak��I�O���(����(0�i>�0؝�\�y��or�.�i��Rm��n�. �;��)��1bXB�hozH/��x�I��o�K:��������Ŵ�*�i��)t���K��|�Q:�"yc='YV�=)�*˘株R�@7���T��n�pA���d���+�d]��@L����]m�Q��A�'yH�%3e+<+�l��y}�5K�!��:��B��{���n�i%��x��B�j^6���S!unASW��<�l��?�Ғm�Ɉ�k0nDԐL�/�7��uHpYCwe�Ǌ}�6�95����D%#V*���|,�/ ՞ �ܭ=YV�:�уʵ��ژ�r���j�Q�>�����t�C�(2�\5��e��C�>����W�Z�U��a �p6V)���!��}�[T��L�˪��KB(� v���]��+G	����o�g�7?�=���.I�9�2���B���=�lq���w��ݞuv������� >�]��<n�ql�tN�0E@��X1Y�[y�DM�-�J�v�t�B ���-2-9߇���̈́\� 4it��J�p�qŮ��&&"����N*������[����)�}�'8��K;�<�-M�\8���uqc��x���O��c6q�����?�Ԉ�-ߴ�MGp�����LY�þ�c��Bd��W3�Ru�F��C��I�t�A&�b�mЩ��ݰ���{��	1�n��ޅ� Ѯ��Yt�B?��a+SB�ǴkQ�@�����O 찖p���2Yd��̰^��4z��ע�Y�(U/����<},�s	Fe6�y��1�u��m[�^�	o�ő�x=�k,WFq�3i��R��2�G��[E�����̢��Y?�်�ںG:jo�ڞ�����sY-�*����,���b��EL#%X3+���U�����l3���w����2I:i�*u;_��K��
?�5*�/����!;Uc�]JQ �(,�I42^S����f`�p�g���D���m��~&�/ƅ<�.�'h����Ǚ\Ì�l�G�8RC)��N��NP2K����ȕt��fB�?�S���ۨ(��YN5�w�=������#O`m)(�w(6C}p&Ѯ_i�=�U�HUfN���[��v��¬G����K���p{]D0Y��q'������i�l�tި�����o01"�v1��moY$.^+�΍|�b]H+ �f�%�G�U��糥J�IA�S+�oC+��ʪB���3r�o��	#8`�M������^��~>IM�����\si,pg϶��W��+�^y�-+/����Ǥ,��V'G�i؎&{{��T��BݛJ���~��r�����&@�5l��kh�#��M��8e�zh)l@���d�����������6Ǽ�ZO�&�}��VV��<�����������*�e�s�0���\ߠ�Y{ju�hٕxc�+�{�J_�L��i�@l2��pKK��7Ý%*�	b��g|KI����R��f�����l6VU)<=�Ϻ��s(j��4	�\o1�$1A�"yőa��d��e�W�?h�b� �R�g�I��8?R��-��2��8x�O
�%��:�q������g��� �� 1����X�hw/��S�{��{��f_w��T+�p��X����К�?&{�@9D��YI㯺!���D~h�.)ɔ����0NJ�uE�g^��&���+h��.d)[��i�fdX��>a�3��ځ�t�ݙ�ue���p���6�Tj�n2�&JZ�IJ�׀|憢�?�ZnD4�s���Y(��O�F`���e�`؃Y
��#��ǅ<<z��?#�b��듞�F����@(�����b�N���T_kE��6��x�X+��G/���파�5�؈R�u�/}W��ZZoW�ȭ�ʪ��jm���$�e��٦�S"��"N.�%�O�϶u�>w$6KSL�L�O���}�0z�>#�Z[5'�< :1�x7�?����8���]]�"+��(�y����u ��9�ڵ�r#?"WL�U�������ީo���^i�"}\�xT�e�Q97R�[$�*�g㌢��K�u$CЍ_����ɢ�us�=à�Gq2��N��d�tyŉu��P�G�y���S��h�Lh�TO���������S�:e�@+�9K���]��Ҳ��gY)���l�������X�i�w�tO�f�'.F��L�쉒}j��i~ĭ�[c�GzrBN:^�� 
��T9�ls��:�zm p���
�Y���u2�^�pqR�7�4u�/T`^���%{�&�	oI��Ҿ���<y�8�8�{j�\d<��G�C�9����S3����&���bv�wÂ�œH���d��qZ,�_�A�x�H�GG@�V&��Ӝ#K��2�N���*ׇ�.�@��*Ἤ�ums�`����kTB�K�U &�ߛ:��l!}� �Pby�9����$Y�_�?�O����7���Ӣ��>�v��w��T\I�-��h����捒��4���*x����B��V�e	��,�O��.n�JAf���l��vs���O`�j�8^T��S�_?�3�`�|��'O��u�@��D��ɨ�;~6T�r�_+���������-��ݐ�8K��H"�\+.e����O��z�^��Y5@<��}�S����l2�w!��?�ȊP�0�-0�6
�\{���~�赵�k��4�p���vtR��l�����:�$��������(�k��c�80���>[G�Kt��vF�T5":�^��	���zF�����2��v::�V����]�\v�(m�zRP���i)�茑������c�*���ͺ��֩T�4�U��pE[�8Bk�Ul�F~~R�W�n"����m"��*��-E�b!吀;����PO����b;�r	�W˄A �M�� �B�9�� w���u!ڱnc�r����
��:����7ۆ�9��`O��6��ַ6�]K$8���j�Z�ʨ���0}��p�y�t�1I�>>H�����)���QO)�&��'��G'@j����X�iX�q�e�%F5�)efy�_l� *UV}�2�����T�.?8�LI��R��߸7\bjx����.�Mwn�� }b�P���9��1��>�:\}_w�8�_��5?��V��ʩ�qU�p������_�aG��*���_w\H��J�Ωw?��E��5i������x%��y��3)9O�,Sb�I�wCt���T".O4t�>|�T���X6R�������`��1��i㝵|�ʁt!�\<���d�X�.o;��
b�k������i��7FZ@O���[��J�����S 3�9P>�P�C	`�k�^���"�߽8�:돕�@�1�FEoM 4�A>i"����j{�ʴ�Q��Yx�o;#c�&��Dl=n�H�K�ߍ�|�h�pw�+Ae[=h��[�h��s�&/^��l&��fm��3����d"�g���q����1�ƔW���R�u����H�Zy`y��`�Zz�%?����Oѝ����F�ݸ�ؙ�5X�Wf$�U�|�����=�}6�����1�*������^6�h^�Q�ָ�%�2���yd]J�K�%�Z���6��`�d�~iZ�-���^���� Іۧ�� !��nG+1$(���!�թ��.6�Z�\��O�wE65�A����&4B�Ԅ�q
��(=Rѿ�%������7^�.b��T��M��R݂��
y��#K�]��[��x�����u���Q	��!���Yx%ӆ�>���U���X�� ���|Wf9Hq�ԵsJ�q!������MJ�>5��EO��ph|�5|ǚ�v�Q��-�0�g"���c��t�9�g�Dc�g=R���jy��wHŭhGQGCt�B��d�	�{}�H�-x.t�dY�{���b�M@����jӈ���kF��.�_�� 3� 6A9IE�G�8>��|�Fו���^��`��@/H�ޔ���Zq�ܖb���1�tJ��k��D.�:���׼K~�%�Ƕj���d&'~��v�ߴ-#��och(����� ��UO��yԑ�ݼ"����6m��|J��=[�Ш�`�Hy:_G�	qa�:3W�kM��n8+(���Xi���� ��v��gc_`-:�� f�h�I��iaO=�P�H8A�$	�B.b�?��%DˇWo���'��J����x��
U�f"��G�hHw	�V@�!�x��Y��xv�2���;�Ky]�������!���⧹�]3��L�C���d��Ϫ�g�MDG���MN �3�7�5MF�Z�݀ŠU�������y�����pH��;�PJ-�ul-�/!�sk���2�4
���G�c�ԁd5�6\���U~�,;���(P橴sU�ۧ�T�.WN	z��B�
t��!��5+���YC�����P��z�qˠ�Ջ ���!���kzƪ�-.���)���i7�4�l[]]�Nc�����N�g9�$��4�\����N�1߰��-�;��N0����h�Q�	�-�h�<���b��;��o�R���������.�%���]�F����B�2/��rd~��I��QU�1v� .6�ːd6Vv�׽�E�&����9�uh��}�?�9���?�3�"g���!Avr��ð;4�m��B?���v���n��Lj��Q��S��}�X�x�ZY+<?r�W��H5�>��?���E��8�v"���a��H�;c=0��Nz�F15J�����1O?�����\d�i��TL?����k8I���_�sj�B��!g\LT��P����ٳĽ4��^>;ޘ�f���.&=w����))��^��!�p�ݮ�l�kG���R�:�aM�^���|�e��9J�8"9�e1���h�D�G��-E���pE�J�g<����<k�02��c�1�3(DbM7�_�=tBs.E�H���
����!3�9lf(X��v4��^{�ڹk��T���۷��ƍp#��K�$Z(q��C��3l��r�崥�8'cS����6��4�0���xB�XiS?F*�%�
 ׆>{��N7kS��aLm�h� ���J��8z�q����l?K2��j�X�7 /����JZ�'c7�JY"�MI���_�ec���n	���#B����$L,�j;��Lfb;�
$?�n�p���]7�b��I�݋ؠ�:� H�w��I���n��$������O���Z�Oyv�p��H)\�f��P�R��kw���m��PŤ]��'TlK��T ��+m"-bшk��V�`1���$��Ĭܡ�eQ�G��GP�˝ð��F��`��)VK�ҁE��O#��t7/�	���k����h%�����Gx{�f�%��˞3y��(��ؕ�rn��\.XO2y�$��7J�K?~9HG�F��AIpz �7݃�k�\�DX�rh}{�Eݜ\V��߆8����?��+�7�ն��G������MX� �'eb�DP,�s��θ.��@4S0
A�v��cl_�z��D�))	���!7��[����A��HpЁ�g	���H�$�"���ٌ��_'���s�|�6��E��:i�s���	��_�K����b8���ؐ�Q�Z9���(N$�=�;�S���Ö��'����p����^�rG�!.����i/mq�j�6sz�#��vX��!�t�8�2���,���XU^rU�}�?�����".	<�4F�m�����'���5?j��/"ق�����ڋS�d!��+ie�+�|�|��aX�0��@����a6~1kp׸��T��IX����zQV�����Yǘ��i�ſʉ��)���(kkn.t�2۸�(C�>iϹ��M����ҿ��M�x�3��]{�%k���n����p�Ң*��UU���1~���TK_�h�c~�as{����H�+-���4�����%���ZEI��b��Cj�����Qbr�736����a(�Y9Т\�ݢ��+����[v��R���v{v��x�l��mk2\9�k�C4P��fw�Kw�V���cJȦɩ���wm�/Q������8a,�@��zx�t�*r?G�L�sZ�	�-S����W���D*�y�1��·A�e��_�Ư�)7��L��~�y�a-�%�/%��$�&s�����P�B��F���o�>�չ	6f!�4f�]ڈ�"�.�G��"�bюD���~�n��^���:��27�{�xM6����"(�ղ�"�.AV1_���z��7&SF��!4{����%L�^�+����дe���v›��{��!2�fJ.!��n��3��uҒ��A��4-���5|�q�,/�l����H��6��,N!�}�G=��D x�8���M�%9կ%=I��|,Dl�VpT\m��r�f�!%"�Sl8�j̙�k�a��ITI��;�f��9 o���N~!m�:f�M�HX2�uzڧ��x��t��x�����A�ͨ7c���e��l��ʛ�C7�+ͩ&����1حX��d6�2CG�mu�T��{s��}BR_���1�)�᠌��(��i̢��ZL���Z�_p�Y�3w/�)K�r�hRg��r���(05}�4_~7ک�Z�V�'�~"$�a�3� i4���0C��aG��V\^f�V�m�Tm���L9��b�E�#a��.Y��[=-���5�
�z�h�~�6��!t ?0/�,//������5�AB�
�J+�N���rw^d���� X���h~�m����\��&�@N1���}a���� ��.P��kC� i�i����ԤZ��̧|�W`"�Jry�
��ǻ!�����10�~S�> :�����xe
�����K�a�Y�C:QĮ[��N&����9�U�� Y���{��N,�C�ⵣ2�{�7F���,u� f��� [�p?	���b��
xJ���%e��9����hv.H�������-[2�+��D���ߥ�<T`Ȯ�i��>p��F��	�p��<$D��J�|�簜|�,L��)�)�(��\��l��OEI��9�EMVY1�(B�&�)�	+�,]�3���4n'����z����R�<���ӡ�6��s���g��q�Қ��Νn�&LS�d��d��!#��&�ܞc����>gւI�AeR��<=X������L�˧�~s��D͈�ل������sI�bi��dpS�֪�J:�ߗ�������7^�t"���W����=��e�9(}�G,b?����hqρ�xgL��YD�H�c3�1����5����`��n"��9� ���c�s�"���m�)g.�4�p��'���L0���]D�.��R��0��5��h�� M<�{�m^��\P\̞7���)'ϻ.����i���܄�k7��؆�3<����u����pj�#R��x"�!7w��rY[!��k\���ni�t3�nfK�
��{'����#1U Hn�?r����H ��WI�*�f�.�7�7x(}�yɮ��!�W��|��a�/B��-ElF��P
<l􏖖��X�j �R��_��U�eJ��wc{��o��k����X��N8�]�m"n����	R�V�%�n�G�J�`n՗� E�d�ߩ�L��6񧜃��i!5w��4��u6�c���Q�6�����,by"��?����%
�:W"��:��gTF�yN��^�0�Q"{�*˟]8^��զe�W�$�9H�v�E���)��c0���r�����eչ��=
\����7�6�P=1C�N��x��O"&$�}x�����VWhCt3d�����U}�Y~B�^K�Q�I��%�N}[��5ߗ��#\a�[x'#볱M�F텷���7	�ɿ�i�]B���  ��յǵ���}}��ߤ[d��Ɂ��8~�s�K#G��Rķ:5[�r��r�c	'UD9}L9Zy�*�y5P�~��2����E��K��~�{�Z�K���!홎o�):ܾ�m������aB{D��?+�B�RB4�*M��sSD0�ة/<LA��'ׅ���r��饌��S:��B?O*�f}L`5V@^�4��d�n�.�����L�Q�l��2痊qO��C�����CKeӳE�A��9r-���d6Pq�}��������t����=��i�2��xE{����ZwR:�6J����6��N��#�/&�,6ȇ%�g���M5���N�����K��C@�I��y��%'L�R\�܍�حX"�8�������J�9����Jb����U�md���lRlN�|������q^�a�X�����#zU�}s�v8�b�RP�2*�����j�Ι��xr��o�Zu�h�= *V㾤��r���G�wL�9qu�u�ӑ:��������"�BX��f�����P9��Ҋ*&�f�R�2�V�p���dѿ��@�'�u�W��ϓ��>Q8Ҁ��z�b�������z�"����W����+� ~��C^��K�M_w݉NN�9��;/Jg֚��/��3��p�JDv)�^�AF���5-��i��*ռ�l�S��.��ԣ�8�َ�Q/V\��̀"8$��{z�0���>����[�iL�"3�ݵ:��0ܵ���SO�b�/&�~i0��R���GZ��`p�m��^j4�/##(4��(�B��Д	�xs�D�M2���9r�Fi��74���%/i+��-ǜ�G���5�p�آ�C0�9$�����w�B�w���}68Z���q5��k�YBC�i�U�����,1�-/3��:�rT���ڈ��%��`i�������H�R����!���]�׊ib�,5	͆2���':]��#5n��,*�Œ8.��̘Ƽ>��#�9�h3���]�x �hB���b��ŉ�h�z�����K�"~�����#"��o�,�C���*����F�C��t^�N������`jX�1�*�M���� ��_�U��Ŕ�juo��������������I��7�0����\��\hIʨ��y�1y�y3�� ���?�-��$���K���!��肨}��z K�������B��y�{f�=+���J�A�C��� �3�7j;�O,O�v����!�d�Ȍ���ȀK��msv��ɌoYc��T-!�t��B*�=�����<�S��?+"s�D��dc���N��D[pt0	%fx- ��5�:�b� �~1?�=7�A��f��>9�S���j�R����0)GuA��8�#�!��*]g.�����ͣ����֠�:��jd�I�|�6+�=exJ�Nr l`���:5rNy:���ejXUҖ�~�`�������J(��(u��|��9N'԰G�Eb�q4�p������ܰ��X�Nl��@���#a���������S�эm`ʂ]�5x���}��lc��2/Bo�
@����ɨ2�T���՚f�:|h�J��]�z>�c�-�9�*���D}1*�%=�d���Gt�`��gc4�D*��kVi�=`�r�N��v�w�����D[��*�^��f,��`BE�	ʎHo|lL�r��CF�#ە�B���u�	�_j�#����6�8���=-��jA��4�wH>o:INq��v����մ5�V<�;J��C6��T�-�!��I�b���l³���>RtXM�w�E���t��c�Ѡ[��C7����kڋ��.�����0��WXI���)��J��7ݳ�)A���4���y:��h�ǹ�D_)p����9����ɻ�$�Yn�w"j��-5�)�����x�]�U癜D~a���
엻 6�UKZ�	�'�g�x��#묇�� :LP��ꩉ:ob~��B�����Z��?w;y^_1MJ�N�L��
=�P4��}��R_��e�[��RD��=n����j�T'a�Z�9�)�����}rO�P��0�9�%�?��_.ہ�gO����R�W�[��샙J����"��8�w; a��Q$�5�sbPWU~��-�#^�-���6�yf?��ۓVS!7%��m�3���m�grnǏ0?d�@:k1�[��Y�qS��񄉟����x/��T4O���Q�|Ԗ�g��s~-��<j����)HR^� �+BG�Bwe!�����xd�������0؛�KZj��=H����T�3�d���%��
P��~�f֦O�gr9ҵ���4��"U��4��ب.\���ɝ���2yg�)]$̈�a�8����x����V��E|�7փ���D�����s�ۅH��uD	R �ȇ�&���:;4x�/L��CHB�.u�C)��J��o�2�,��}���h��էL�"����n�bFK����Ɖ���Xre��T�`F��n"������Z������o��t�9M�-<MWl�������[�w2�������'<����%#=����C�v���b�P���!g��b�FI���d+1DYt�O��/,[�#�����nܝ����d�[��Rh!�S�Cf�����j���W/i��%��b�C����}c�$�.�2��6^�5����3��z�"���]�
�K!�1���.�z�{e��`6_!��hdm.ě��p��gn��(�n@V�h�p�y��>�
���ޛW4o4�z
&�5�Y��W�(WJ\[�u~�5LN�ai��UudIjX�
�ǻ���v���P$LJG�'a���e����K9~��׌���/�lb��Qδ�����=��a���Q9�ca�Zi^���#ۃ�Gx��[)�o5���H�������^���Q$��LP�{���O�w���q���WB���̄��e=�g�"u��5t��0�Sb��fOJ׈�U��FK�n^eti�>q¬�W��I��o\�����hr�<x�7�:�<{�'a�E�L	rD!L+��5w��Y#I�� y�Q�3���jy��'9���LSE/���%��� 2��Y���V�Z�Jw�%< ,�~�S͌���������%��ZRG�܌�Km3$��a"3��$���۳`/`5�@��b_"����n��}��C1�]2^;�}�$���m��������u���u��W�/������۶5����-�>����Y8n�Zn���p7/�WX� �@������\/ʑ�BD�x�[?O�p���iE1u�ٵ��)^L'A���)g�%c��4a������ZW��y��:�u}�@]�}W����O�ħ�$i>
;�Zc|�>ژ�[)�����K̭b�L��r�2eB��&��Q�b� �B��N, ��A�蟛M\֎���[�`�i�r.���ܯ��Pha�K�������=�F�~+&
lP�N����vT���-x�������uI_�xt�,�'��y�@���j@2���E�P;3���H�=%b0�^c�
�&��-����G�k�����a�˶��:*�IԴ(�8���C�9ϫ!g��7�:-��aOb8��"\���nr~.ܛ衲IuI�����Q=1r�������<������0���[�[�]��c����v�X��K��{l#�E&�0jE�Q�?���/��Cry���{
/Bq�=���Ն�_����f3��J,C�;^|�v�If�Lpu���Z� ��c�p����S�X���O�(�:�����J"�o
�)��M{_����7�E0u�lZ�w&�h�8�8hv����ߒ�kWuZdV�s��(�_ë� %ƽ*���9��(y�q�x�l����2����1��3���	��'��x��]^�_k'���:>�.�\�k�A�Yv�"�S���aڈ�o?z`��S{�N��Ju긧��O��X�9aV����Z��:�~�U�*����U8��?2�|���k��^��[�z(x�y��byM����;��P�"�0(��lO���m�ti��c���z�����L���<�8˒�3$[,ʣ�2��:|�#�>W*$����Ŀ��v�(�Bܡm0�7��{�s�/uC�-����)c>�=���R�`F��@�����\���>��Ԭ�J�K�um{��QX���g&*.�]c�jI�tt�8A��8���/P�����o6�p�˃9>s��L����,�Z�*F,���ڌG{�'�C���z�����=�p%Q�5��q���{�$����\JoJ���O��'�-���G��΀b��-oa�{�oeE�~�i�!�	�������#�����(���H��.4aDbck�R4R�K���X�{�n�(�ϕ��j0'�T$J�:�'�bRZ+��G�@S|	'���/%��-	ӭ�Ȉceݏ�;:X ��WjMil��Z�?���=�q-ƃcK�M�=���B� 0����w���]dq���7�3���@�[C��o[� ����bՙ:���]�2Nr��w^�S�����8LyQ��)ъC(��f��dŒ9�h0�l����Z:[�WJ�u�Qʵy�z��o`8+��y��&�~繲�(	�֩y�:AR3y��d!�[ˣ�U �n��J��D�2����^ u�J7����H|{���@t����>t�k�+�|�9w�TW���Prou��_��sw��z�����6%e\4&~��#��Px޶���U���(�!�����3 b�CL���WJ���:���SH�������b���N��J�b:Z�;t8\����Z�(����	*0���H��d}Ƚ0�Ʃ`�gz�`���L5�~+n�.���MA{��,+��9�vc�Y����׬튎�y5f���3�A�Y�:{A�L2~٬�p۟��MX&eR��y���G�k��z ���O#ti�b���Qn�w$_�~�aA�UH~�F�HN�����Mw�U���������f����j�۷ץ����s�2S]�R�X��h��n��x�]$�\ J3I�G/�Wdb���x���L�2�`!�h�(��ɭ����&��-�p���r��qN|v����^ܤ��t�&1^�b���m��_V\�ݽ�$��Z��[+�ZKvaHe�l����?� %�uז;,p��1n�Iu�G)=6���b����?B�u��9�<������:�A��f��YՏmB3F�Y)�?��*�)�JA�~�=�t��$��YԲi��R	4DźA���n���\��;3��B��U��8hxE.���ڞ5<��
�Ǻ���=UK8��*�:�c\�b�!1��S�A�.��N�`�,Q=�7�U!�L���ʛ�L �]�n��}2���w��~��g��]�U�(i��S��,͎���Z��$/g����%+{�šM�+p�[8�x�"N�x�$H(��,���FH*t��|���&ډ(�+��;�jU���0�4��R����a���P��M8θX�SJ-�߈�{i8��M� X���8$��J|�B��ͪ���94��E��8J�Z�gݞPK%eٗ�S��N9᭗B�X��YS:�B������@����e e�Ǜ�
�(�Sҷ��[��17g$��*i���0g�.cW��3����e��d�-�ٙPʐ���2�|��<ʪ���@���r|1��3�5��p�����`���3�{$�K�,�|�)X��V��C�P�ڜ)P�0��`�]]^}��!\�m�:���$�m��2�j�7� Ƽ�k�v 3�~�]���X[�UZ�������5�^C��}G�;%���k̀MJ9��F�R�28��0I�T�l�0�J�\���:���x/�f/��E��+�Mw�\U�&$��T	�ZO���b��5����n�=�+X���,d�K�qe��[��N�pM��r�Պ8�e���)D,���%d���a�RK��SP�L�%�ư�}�Q#&�΂K�u>�P��tj���^�Q,��2|�+��䳏�r�0�2�n;�����% �E�M��Ȅ����t����2�)�,��W�w�~jL��<���T��]'�	���6���e��c9�|mI{>���ߜ^s���.�$�(l��}��FEWU�>.X�5u�������񛢰�.����ٰ�=V���M�(<��`K����V���k���.���Ij���Wەg�>���8E^�߮��݊D�6"*詡]QQ�Z׃��y�V/�X�'$|y�
�ɟp�]���!�5P��ˉ����O����&�u��P�S�W�~մ_z�*���ϸM�Yz��_�+��oϢ��	��Q��=Gǲ~��N-1��|���~&���N��8
���n�#,����,��k� �5��qr�U��D#��P+`���7>t�N�K�Kl�<mm��'f��M\����'����풼 R��J�۫�W�Ϫ�3$˱�5��w�f$�&�^Jʈ�I�c��Wu��e	�[�1�1��0��m�í�ȵbJ�yPH(��CrsޡV ��ok22Fb
t����;Щ�O<ѵ�NH�H�`b5�d��s������ғo}��j��9��+�D�4>P5A,A+�|;ė}���qt�a��K>� '�4I��5ά� �(�b�Şb����B6��-����Q�)b��=�k[�9��!��w�B���F�༧r"�UT��'o�[����V4� 
����nʯ���K}���a�"xvL������`�݆V~V�HX�$���<�Az0�;��KM�7��~���KJ���	NQ������C��Q?�-a�|���_$Yo'�����ev���K�zu���U�"uk��]�#$�LU{2�K~*"d�������8Ǘ�����g YQ�On!�{��E%�����I�`�|���Ź�ō����׮�g�ζ=�\{|��S/,p��Kq���g|K��(�e����~�FR�:y�F�$�Dd����"�X��|~K?1AJ-k�~�X�g^W�1�O'%�I�J��Sx�r�a=���0&�M�����ċ�i!S&�ޏ�͇���k�i�)�%&�-{7���B�����cG4W%���c�&p�R���+��T� �!^ѾGXy^�3đ���h�K��l��fGBo�م_�k�` �V��q��x��r��~C:]I�8~e��G�"��LI�#˪>��� C��!�yy;��4�.9�$n�<�{�O�Y���*"U2��-�?��j���-!ւ�Y��F���?��:��2�!��3ŖVʈ��?�p�<m+���9�6���M��e�KP�h��q��u��*�Q-��,o�۽�6�]Ӳ̪߬H�t�4��[�}�G$!��Ǎ�W��UXiS�w\`�_���J`�s%���Q��'
�Mg��1#��V�_T�$�J���0Dos?����)}�YÂ���(ZM� gR\��m��y/�Z-�a\^�hg]H�Xǭ ����ɞ��)!z�;v�,����t|3��C��qCj"��'�y؊�,��׊z�X"�G^��b�7�������$��֗~��i\h��2�,�</ϮY�~V=e]��)��P�k=�a�X[��6�G@��]�o�	�`UKD�P���F��ZX�b-$�xN*�J�詤@�r�C� ���z�8�Ag��~��d�קܖHy���u�M��0��)���ye#x��a7y�n���j�3���z;����a����~�|j
t;� ��X��#
Om��h�D�6�;K�Q�S5Z��'�~Ml(G��8�p�����5��\UC��w�?Ș�1�:�"�5Em�����Y
��ix4"6��$FV&�j�H&�a��%A�/G��}�ǅ'4A�:7��0.�I�Y6�͍�E���&0俩���i�:`=mg�˪�s[wG��Ԛ�:=O���,���M����|��?^����*��٦��r�V@�Cե�g�� �P�h�tf9Mל���X�P�Y#�5����ݷ@˹��Vl3��s�V�2@����_����ttC�,�� ��u��O~�$|��?3��J��ƀ����E�2/��Y�ia�Q�*�c?��y�7�</�f*.&��f��L@\Q�CcU��G�埠,(`��bBc����	L��l��n���ū���=�ac��^��	�-����I�뚿�B��Q��lY�'��!�t��5)H]�\��+� 2���ި<�_��4i��b�����7j6Bn�KT�;����v��)1���I�����>�e�ѩ�w�y=�~����;�E)��
?(=���d`[�;eN@�Z��Ъ@�9~���c`�A\i�]��-���2܂ݪ;vƯ��0�^�ɒH��%��[N�ˮ�H&���9f�n�}H��$\���O��=VػFC�Z��nI�ߪ�Y0�/��e���k���Ҿ�^��8�0�/��-���|���Rde���^Nؼ�'e�l�\��E����AI���Ո����H�G������������*�g&���);��!�I�3	\�B�7#��,���(®�Ge���h�"��W�/�S�u*8�<�+�$<�ݣ�܆3六X�`K����U,�:f����Q/�4~6�]�����Ѝ��A	W������Y���%����F����Axwh��p��ǟs~{��:b�ڴܔ�C�*`�nA:�{;K*Ҋ�Y[T��u�<w���_���<��V��M��?�Z���m�c��* �[ip�s�Soq`�Ʊ�e���7��F^L;3�@K�(�y���7��0<�Ti�Xk&���O®�-�6-�ÀEB7_|�
�����2ݝ�g[�>�>T���2�k��|m�m�UG����z�%�#n�6�`&i2��-wawVb� ���=iw�;��\�Z�s�ֽ[+�;���Wj�b�a�2�͋�q��6+�A{ A}�\)V1��Cw���-�M4�ݛp �1��lj��n��$�C*%������4o�ʜ��ዖJ]u��?���4b��x�C���u�3<�N�m�[�k��=+�R�s��4�v��X������۫uW����T���s����*ߝ	L��M���%��`㟛��N�*l��CCj�n�o����������	��J����n��_���`Oh���c兤��t�5e�>g;P(�E�}��z�Pg:�YGtDX�E���@Ph�l[^;���a��A��;?|�;$���B�6� 2Ij=�e��m=� \~��=wvLc`I�V���I�aG{�T�,��)�{U�"8����k qu~�$֤��Ծ�*/O틁�����ƚC���}�ji=��jJ���m�\�5Hm1��v'���c��$�'5�~;��B��PN��[0�,he"Z!E����͘�F�ş��g�Y���ڣߚW����kϏ����ڐ��~(S��y�Ì��7r�D!���AQ%����h�hc��6�tto�Ui]h=z�\���s>��o�Wx<�W�s�c�ۭ����5g#�3z�C�nO�[Tu�}�i����u���v��r]
����]\�[�J�0�����j%�8���� �B)��'Mo_��=	��?DW�)Y�r0�ד����Oٴu�`�.���r��tj�L����LMa�(���ԚLƑ\ǹ� �&]2���R�5�e ;n�M�L��N����1o�r �O۞��@�oD,aI��msiP�;�Xﵱg{,>J�Yj�ۅ�औ�B�8�3U*B���kDu�%h��$)�[	#�%]�3S���iK�\��V�%>�
ή�P��wc����WKd���.˺q��(�_�JgD�!XR���o�hIx1�4��U:���?
�t(�������NYS���	�����"���"FbL�6C�FG�\8Ix���~���~9ͯ�ʶ��U��cn\�x���_��<T��a���^l�W��L�*�w�ݻ��AG��!F�D�PJ��΢fA�4�x��7|px`�#�@�S�$:�i���:uJf�z"oH�X�"�N&_�=���4T����D���(��O��s�;Q�_,!��j�Y��p�IF�2q�(��N���4�ȩ7��9W���������3�y��#���o�.��5-�K�N�u�d���&��D��=t�X��J�����5�vBr��IS����c�����,5�����릣Q������u^���ۇ����g�-�a�f{��W\��	��ɁDg���)��V���KH��wi�D?G��;FT�<�<�k��فt��0'zp���DI�%!D�<Z^�W/f#M5��d�^c2Wf ��!!�M���Q����δ����M
�4��vߓ�]pݎ~�Q1M��ܥ��C���R�s�n���P�3�3����?���-�$ l0�PA���]��~.��OrGs����q��7��ȵ[WS���4G���X*ڭQ��f�?]�ae�?aP�*�h� �Xn�D�%��������~eʾPn�+���p�@p�t�>J��7ޚ�ۑ�d�N�j�5��HtJ��8e�:`���%��r�52d��x����kΧ�߅*"��g�_0���^�h���g��Ӆ-z�O�p!�1m�"����;8
u�g}�Q���w���k�_��`c�'.`Z�h�����[�q��e�!�����E
�3�.9i1c0^9��%���"y�(���-��-�κx�h�1#�H��*:����3��r+x��X�X��no����~2{;�T���C+�0��&�P�a�|�>+h�p� 4�y?b��c,V�i���#JR�g"��%V���ca���-W��+B���G��0����A�K8k)+�ŋ5�_�hʙ�C�
�ݚ���ࢴ\��n���z�X�;� 8� ���@��#"��<N���VV��0�t��`(n��(���nF�;��t,\A�~���O���<tű�1�f��|5�~7������Q ���t\Q2�ջ�\y��s�a���	�7�� �U�~$�O��#1�;K��K��A�H�O*k��;z��Z��*q(R�[���̣w}�K*f'a���,���ӱ��9�Q6�C뇭�����P ���eϻ�ë%��gDcm=k�f.sfE�8
I�߿�X�$j>u����5P��ey�X��#�T��U{e�
��hR��}�����{8�m�Qc�'�;���`��ޖ���ʁ ZO"�Ȃ6P������9�6D���\��<���`B?,��g���&�(�Pg!�/�xm�#��A�e��:gcE�k k�;}*�5�$pB���ʝJ�ŵ���^u,?ۇ��ݮG_�y5MGG�	O.I�^�[D7a������{�^����'�г��ք�R�X�0�Pﴩ���{�DM�H�uζ׿���+��`_��o�x.�?����H�~��%ց���T�V��+��6�8�ϛ��I�/6fg@lkwYO�	�!:�r���0A>�C�b0ϙ�z���>-ohޛŨ\B�R���[�l�q!��p(�d�h����b���/n`�r]B7��������V�P��T� {/:�ED�H2����<���'�v�]�]�ߧ�h�5W�w��$��'BB���wV	Ztb�V�?-��,"��sBT�P(�����Ɔ�f#���TȐ��{��2ۊ�[XET]���H,j���i�7/7}Fl��"�^E�	h����'%�����k{l�"f�:f"�ɓ!K�v0������B޳hw�L���@���V���I-M�����)���[��I^���<E�����1��&����k�!L���p�0��uHcx/Ѿ˹]�sw a�#9�1��|��	y���b��OJ�!ë���-œ+i�u�w;��nJ�҄�:�(��|�*�џ��g
��4ͫ�����%�f6�\j����R`�����1�:�9��?�-����d
���׭�1��=L�mx��9�� *��#\�?�;t��lN3���3��R�&��w+�(�bkMe� ��%�4�B�o�42^6�t��p ��k�e��hrAb�<֊����e��rړ)����Ċ����l5�[���pf{v��Xp��Ѥߎ���IC�o+G�����gE��b� �}V���g`,&��W����g�ʊ�W��2l�)���m'�8��DM�I<�I�.��R^��s��܈R{٠p�ؕ�&q[_1��$�{s�7����%"��`�m�aT9
O���~-��v���iR˭z;)�N0��
wB�v�<n�!u�b$c�ң!�z����fN�"b�Q�!�H��J\M��Ų҉�pQ���}%w;���]�X����
��R?V�Ed��u`�Dz�YG$!�6�mї���n�*#�����Ӣ��
 R�Q�	X�ɔ����&)B�����6W���i}�����]��J�1>IL�d20�Ӊ�X]"��2O͇ ����R�D�U�4����U�)��t���טb ��64nZ�a��E�Q�~�辈^�A�����  ��Ty�+XM��Vk!�n��ԼZ�ܕ�L��+kI���OR�0"@�ArOE]s�=���?�A	��U����]���m'�Ή�Qj�un?fêO�Oy�+�bgb��X�n���C�h�M��v��mH�Q�؇�!������2���ع�@�0J�A��Ek����擜�*�!���1�">��R�B��,���-����
�7����O��R*��y�}�	�1Gnn���és#���2�A8�	�$.�0(��'6T/���K>v\�}!���?L��}�|���T%�}���-M3�6�A����*`I&�Ғ��$f�֫��_���{�NR,��ɀ��8�ʧP����0$��lt5ȅm̬�gmq�b9|�#�W������,���6
[9������I�Vh���� I!*�3 e�	��4��W�����4�/V�5��2u;7*��c$M����,��"�v�5��L��_T޾��z�[�*6>�����"���#��$�K���P��J8�x[Ɍ��j��,�aY�5��{K�K�.:\`3RE ��D�ݪ���ϑ��{�'��B}4F<s�o-m[�o��@�"�)�vȼY�����A���qF�3�9%��xn'��8=(���FN�Ćh_�~4փǲ���>N4���<�4bY�[��٠C�C��ݔl奞�B�Z%ƒ�v�A����ZO$����T�G����tl���>���@����P<J��0f� �	�I��M_߇��W$9�$�����[�Р�0����\\�")g~��HT�2���,�f����5\�y�a����hO��;f��R%x߂;:���=����!��@�>�o>��mAC�n����$���U�;�����=]���<� a�8ɮ���5��mZ$T.	�@Bk�������t�u������щӋ���j�`�<�QRR�9�P�w��2K95H)���g����~��A�������xۭ�K��)��b��r�'?��Xs+��~Ɖ%sl�s�H� :ZЌ�n����U$yӱ�!��A	��&3���#���<gc��Z��gp�f@h���"�5�ä�_���C����������q��M><�*J��-��T�RV��t��34D�)�N^c
�ׇ��R��ő���8�>����z���MNl��,~e��X����%��T�H���Nk���/�}P�
��������gZ���D�#��D�y_Z�"��>�o�� �j�8��Q-wm\��9ɞo3�����:~���r'J��eN��2ڷ�u���,?�x��|*�8�Q_f��P���27�VA*��Щm�-Kk}^�C�C�㺹����9�O2{�Y��ٚ)���+�8�BH����ŀ\�1r�����ϺG/u�����vFF&��;�o�Ab�����#����uO������W��X�]1�p�Z�-�ܵ����R�0����0��+��x7�>��װ�q�r�]9��Iuq�`�GX�����;	TW��J���YbmqO�z==����:�m��e����Q��3���q+����t���0��b�u6�J�����Y�̳��h��B�ez�*ElcZ�P��) �,P�:�z�w�גϕ������6��Jd;���wͲ+(�V[�Yv��H����3���,����8���sX]�I-�S���.�w�>|΃�n~���`4���P�Q���%F)���[�f�x����l�HTE��ρ� .d
��),��7�Ѡ	�EE^7����6�$� �AM9���ִ�ѿڣ?�$�Ub�{�Q{�r�/��+3�8ſ@�K��h��'�'�n��΁����%%'W� ���H_A\M����tC�j�a�U챠	�e���bg0M�R��M��I�P�0�1F��7	�tC˨�8�V2��*�C$.��L��."OC� F�8��F�g�6�ͧށ#]y�ч�-R���X�sZI$֡��?�֗=���D[mן�qX�~�؍��H�]�]� ��ɟ.�m���� �D1s�~��&`����PSV�3{����x4��g�����O|����"̐���\��kܦ\��z��|b YdbSj�GH �P+�F�x�-�F�'�?����;��3�K4-~)����\=���A|e@+h? �]������:
å��.�s�U���C�ҭ���6�>N�����y�=W�A`�˫1��Ǹ�ͅ^#��J3hT��An��h�P��>-��߯�p� �t�	u@�s�X��%w��(�#�O���r���.�"�|�~��4f���cu���i�*�z��KKNm�l(.Z\Ƿ0Q1�f��Xf�ѥ\�Ɏ5ʏM��."W\N��U�[��q���$�K��.�?�����P�w��i���{��3�.�ؙ�W�����w%��a]�IC��'K��kP���7��.p[F�[��3�fO��7��'x�]�Ź+}����x��S*�����.©}��njZLE.�*\�(��>�y.}���n�^���"X���X8T�E	�RĀa?��1�B�M���\E����_VMJ ٲY;��[3��pd͟నd^Zb��'<}���	��;�[��iK���v�c��պ�a�i��8�F�=���X����&�����Ò��a��M�r�ho���vf I�w
[("�|3��η�了��%�� ����5˞n�^�W�Q$��4��41�Z�h,&f���Z�e�֬z�a����[wҝ.K<���x%��D:�yi�+��n3�����Ω3�[��a#w��ƽ?��8�mQ�[-K���D��<k�_+��D�\���z��aُúo�z�Ѳc�,g������t�a$]��H� ���]�XSkӬ�׉����fx�If�i��aΦ��t���^�H�IԱ�j4}�� o"�Ԩ�Z�6	��U�$.���)��I{Ɠ^YS��̸���6'`���.r�va�b�$�ii��k�Ml<���ȶFr�5���R�6h��VMQm�4oS�tqkEDẲ?Π�g��n���d��Y��;G�1���Q�Y�Y�%��q��X���QU��psH�f`
��sl�fPC���S
�Y��v�]D��q01�3G	3�%���/d�|�a!�}�g���\m�6mi��7��'ϊq_F*�B9%L(�9I/j�2Y� o�������y��ߪ�$�1
����&��T�8W���̲��ٿ�S�;�&n�\ov~w^�*ۇ��h������n���K��V3W��͔r��y*�eD�$���Y�6��zQtoR[F�,;ϒ�l�S4��˪]U&�FB�sFՓd~�y����H�l�r�>*�%��In�F�7ӨM���T�?֮���*?{����QMp@�,�޸���~���'��zT�<h�(�5��Lp���OF=�*Du&�ϝ'Z�ڴ��Vl�1��$�=�M:0��{������p�5~f����H퓼��"�7�M�6[^�t4��3[�����8uS�.>�ł毡�4܅���w�m&��Q(�Ѕ�vf�CM(!O�_�C믿;�A���#��߃��{��v#mM{�yy�伩B�=�zQ�qJ3^:c��Ww�kZ1?/^_����IZKtw?_�&���s�]@Wp�<��W#�d���HO�Y��NFx��	�*ޗ%	���Z�b��S�|�#*v��p�ƈ2�|���u\u�8��CFVď]!����ʤ��_w�Ų6�+�5�׳z3X혚��3��\�Ӛs�!v=��4ĵ;ڪ�r�����8bw\'b��Zн��ƚ=�7���AU�6\7������+ۮ��\���P���|pه�{d��?uXO���X`����J��Jy�g<*�y��w1y�`澒�^��`?ի��M��R��+6�p���� �Y��@A5�4v��΂Eq�B1��%*���[��
�y��dAF���P�*�l/�k7��Rፐ4��2^�L\~�WF]��fC��@DgR�ep�q��r;!`�c��Kÿ��2��6i&C���a�c��0���b���K9��:|^��|�h�G�{�#�E#����T{�D��zc�+d�6�������v�$� ��!%'7J�AD��>�/ɻ8����P���-�Ȩ��M.kߠt�_��$�{Pf�J�i��DUu$ǚ�1v2���Ǩ�d�x�)�_�������63�SYd>8]sD�t��5� A]aJ7}�s�H'GC�h�l�R��q�sK�Hԣ:��b`sg�2#R�g�����?HG
�j��rw��p�J����v2l��@���ߑ�9�X�"d��Ӽ>���t�^��W:Wj�`R6+�\ԍ���]Zz�t<����ǽ��:N��1���/��KvX=^�Fa?5��zyk>R�Ѧ�-yrPN6����ѿ��w�l�Nk&��}v�4�K�D�X�j�i û�
�U� TFzЧd盈���{Rf3
�8�@����k����	�m���M�29QY�ؠ��-6�V���3�C!����/��Qf��]A�/�8�������Y�&����2y0�AA���#󦔮��c��MK��9�t`��.�ǫ<�R\�t��n�$�U�I���8����˲3����U��&kdCmSlZ^�b߹C�n�Ö?h���.�6���.;���u�.��Ģ����i#I=8B�h�M9D������&
�3�q�"��-Cy�T�p��P�լA�[7�����x�N�_�T�k�P�I����#�%8�(1و{��#��ާF�ݠ�������3F�l���>�GW=�tR��o�`jKu�i�0�-mt1� �@��Q�(�l�>G�]������;�i'��|��=�Ǣ+?�����pR�d�}���VN�n��%Α�d��Xb�T*x�r��j�(㌕^����I;�dd��; �0�ٱ5�H���/E5w=��z��n~�fI���pU�u����:ܮ�S渪���y�g��R��޺��S�b�����:�,\���I���n����}c.]_,Y�����ާc�ɳm	��܊y�B�o�ꖞ��!�T^�"+JO�{���a�-��,vyxo�cH���	*b!��]�^6iB��Ж������ј��.�����m/�X�O�\�w�E���@�6R�U��-]\Z�V8hA}]5͘.��7���8�y����:�h�v�h[��\EI^9(���+"�-���SU�zODpaa���T,��tnO�2�~y�&q��y��(�/��ٵ���������ɒ-�Td}�zP�E��������%�p�ɹ�W��LJxAp]q�5�����X?��C�S����"J:���yZ�7��M�{s5@H4)�_�x����梢�+@u���7	�ԯ�ҹ�Bh!��6���U����W�yO���`]Bʅ��R�~�qE/t�ڥ��p�Ǥ�[�'�%�z�o/j�`��� ��+�Jr�!�f��ki;ԯNCv0�Q��0B*�GH�����o�	�y<��_A@����+�T9!a �T��<rV��{^^�c�������4���"�p�ԭq�[��;r�Qm:M�楘_�$;ʆdXD��Fp,=���4����xf"�]$7��+R�u���7���������f�v� �:Z�����]j'����?������K?F�Sl��{���'�r�E�R�tqO`b ���۸t�Y]`�]��`bq���4��0L�b�r�F�n �A��p7�����Lz�À9�E+�#1C���k��U&�]�]�xI�����h&P]��t��p���~L�c�-��B߶9���cjsu��s|�_EstA!��w�'��܉���N�-�+K���+���'<U#�1T�@��:hr��#t>X�!0�ŀ��ܳƲo΃��o,O���m�+x��0[����i�4��Q�XC�A����Ϳ��?{�EƜ=�Y%�Ԑ����h+ �?����#Y̺�Z�;��0��b()54'S.U,]8�o3�#�wg�V�{���r��a�i�9Q.o����+C�������s<<ʨA�;�7���[�Z�Xh�u�y��͒�>��;D�ک�/�z�R�Z>������s%K֏f�>2�V��� �m<nk���'�H�����<,�CE�3|c�"!P.�ȏ��Nn�[��\1����e1�o+���^���J_�?�������+��@x��_q \��C���~b|�ǁWO%���>��}?�
��S���5
�t��UO�	(����)����X�x������%^;P�1C*��CaS���| ��"BLg*<�@�������A�e{%�W�9�e�R�(�[؛b�['�����Eb-WD�����;���V���C��p$�#O{&�0R�BK�Hq�fwY��R��B�<\[AM�yg�
Gx��J�� z��Tu#�M>����2֖�_��Pзh۫3�q:�����qi �A�j�}�����
$��߾��"+eq�A;�9���M�j�LTT�p7��Ͻ��˩�0QC�^��JN�C
�җu�� h��N&�ѣh�)�ձ9�2��G�|�"O#�X��djc;�u �^���nU�:)��&K�ݟ�u�e�M�[��L�`>Y��0<���~��kW
�5G�q,�$�`-�.l�i�,�#�{�J4v���]_�T��<�'�ѭ1�U��ć���ߐ�c��2n����o0~�	�խ�p_���VH�ء�[��\$�Ee���jW�NWåh1���G����*��M��t�đ��D����	��$_ʗ�|��dD��{dŃ�� ��1|�yZHQ��n����ed3���%`�y7c$`>�2Ml��D�Ød{�����D��&��qR�����-V�E��9I:5]���{�I艚�jZ:]J�����?�.v\��Z{�Ac�Y�oҫ� ��H��q�-wyR�� ��HI������}O�|�+���""c���n�s嚂���٧�#O�Ӎ�R���������cur�i%>t?q��y��1F����e�i��ڮ��g4_�v�jc(>�P��7��J��@Ü��re��(���W#b�:�#��/��.s�vֹ��*lQ��;	�6���-8R`��Py���s��?�S��pBI�0�\qbj��3X�37$u��$w�AC(s�)p5�` ��cp�U�t���q��E;fx���m�A6)�]������S�s4�Dx��#7!b����@���+u�����2<��8H<���ɲ��SgFv'qq�9�������ncG�(�B�M�� q<������>��"h��d-��8�%�L�y��f��ݞ��<�]�M�~4�)mgT�H��mJ����UT����cvN/<���9�s���u�u!6�*�ԣ��{qu�2��3K;�1t5�F�F�j�:"��3Q`=E�Y����)9wbF�>��=���d�WpH��!����N�O	a�7dAv��b�O�8�.@K#7�N� ��C6���҆9�"�����1�0���a�{�?�l�0a.$�_�d��p�g7�p�%M{d�S���=ʈ�j���#J��{��=V�ZVo8;b�"p������=SSg��s���j�)�Ir��w$Sg�%��r�/�Z�O P���=w�G�G���s5ߏ�ym���^p�0ҿ+�<�ju�%�v�L�SZ7^�`�<a�*��E��5�Hn���onV��Lϱd������	���� �7:^����)�{)[�$�|"�A��IB�%i<h=迄Q@#P�~>�������"��5Y�yj��-��f��.�%�������d��t���J���^��E=��fG�,��Ë@[���Rz;O�D`�Ed�GY(���;�'�����BhV�U�OѸG�2��X@q������)!i筻�Ξcrm�����u�"�.�Ht.�����|�E����D���Hx��ty��9�m�[��)���qX����}�Ig]�7e���%1F�;��*P%n��ܝ�5v��H(9@��BF�Q�Z�5-6ͮ�}>�abB��b�G~j�&��EwE�z�+6�XT�E�!�I=��)ah%}���V�
FY;����!���5�߻m�I<m�r5������C?���甐I�9v �x���l�0�8>b��7%�l�������p�KLL�g7}�rcu��#٤D�z<�\�y_x^}�\c3H}j)�y]�u�\��Ŀ�gDu3����P�V/�Hڧ�A3��%R����e�03rw�ܤnYwߨ�N*����*�{Y��Kd)L3�,f7��f� ��Q1Y��%ǀ8)Q[�Kw5��A���Q�:#���)C
��7�T ���ki�ӆ��cC�:�R�T6.�Z-�,�MHc�����ݬ8��������(]6���`>���j����n��~X�E��hz��j������I�T�ϕY���Y�޻�7_%�=|?�U��3e��/�`�Rr�G�����jĦ&��ǤK��4�����%Bҹkm���S#�+�b�a�e����v�w�<W� ֐<�g��0Ag��<_���I	]*��G�����w��Ɛ��Czx"W��'��GH ��Ȕ�}L�Լo�=kz7�����L��zGMY�����=�EV �
��8X��y��� �[�暈����k�r����}���7��ȁ��FP0�qѼ���BG�ץ3 �a���ꨦ`���|�X쾙�H�����tJE�52�kJ�m�휧�)!F�综ݳ�&F�i����nWC�ǂm�d��_#Xt�+��O��_�lg�\�;�뜸�H����Ak*�3^wY�q�J]�m�F���|�?�h/�+;wD׷����W̓i|��ɂ񲡅�ฬ�=��(�q�/f�z̈́) XJ�	j��Ơ���^˚
�ň,��2�J6%L5X�x�|P�Z�N�p`Qyo�<���Q���okq�P�D��9�"=q��jE�9�J,��M��}~�L�+X;��d}���v�^��jD�HT�ڔe��^�8I���	�F��_;@}7	�B0�7�ص
Ѐc��]'����9�J=�]��H7;|F��.aS�wo���&xD6��c����
����NO����XS�!Y�ýBu��<!�v{	���%L|wrc�� �M�Y�B!�2�bo��{�\�K���Ou��ȶ��M1�5OQ{7{a�X#-tG���V��t��w����
��׆���Ia?q�G��\��w����T���q���m7�2����{���(y�LcB�E3��Gf����9b�ł鷙����9g��${V�!nY`a���M����'�
���^|�㵙�6`�=��٪�/M$�7=y	��2?E%/L�e
[�N�7^[6{'����Z-��S��l8u^�2\���b?��-ֳ%�C!z�:������?���{�'P�6m�-MѼk�E�N�R�R}(�2~P�pK`�/9�ulLp���zq�h#�Caoz�qإ����<���y"]��̫C��z��dɫ���N����&g� s�~����9M��ةY�^�/mu�Cw�f��)}����O|]���A= �p�U߈�]�!���d|2W�q�����k��Ý ���Aa�[���ҫ���/л���Z�@}�W��	'%.G�RtY�Cu�T=�p�J'rN;~�I����~����f��v��-Ǻ��u�tL^����{4��S�[y��o�n����]�}�m(/n�b_�t��N��#��>����U[h�^���M���b�w�Uۦ�4]#!*u�q��a���}�۱��ܮ��^i&=;?��U?M�#����$x)$F��j�P�����$�C��A{�u҃�J�T{mA	W_(w6*��0q���)p��Y�r��I�jZ���X�uв�s���-���N���uE5��fI��4xWɕ�2��~��v@��'Hx3���cl�x���6�,̻�0�D����3�}m�;��q'<�S7"���k�u@���y��i�j�;r�����߇W�"!AV�l�4����<Ry|KI�"E8��)�0���B3pd�p?�F�X$�J[�`�*�L�t�ޫ�nw�=]�F�\һ�o���
��5l�#��aQ�-kz�6����e� vc1�����p
�=�G,�+`�Z�^�E^]ԛ �q�iv9��q�_�G0Q�le���Ѭ�G��}cq��:qy$B�5s�K��z�/o�yT��Bi��Ρ�'��G��t��DI�x�-`�,���*�w�)�~�|[V;y!/���a�S��}z�u�P�*l�AqM�ߚ��<�&i��ZĮ4H�m|��Cˑe��rnŜ��3�h+��e���M'.@/f�~�c)sJG�&8�6B(��4"SA�&̾Sb����H��|�Y��mO��S &�M�	 w�}O� R�  ��Y��_~�/��\E ڣt�I ��l���W��ڹ��9����d���w��*
�
z��n����畽��eң�1f�0��Ж�8��i2��� x �j+��;�w=��V$�<Bd�� j��ŗM!1�!���F2iKws�����Y��	�ߢ�����>�w�W��$�x��P��B}��N��ǡ��k$ś��Tu�7b����zI�_h�i�X�ڔ�e�q+%<<��y�Ʊ��#y]<�@$d� >l�����0*�H�4.|PK�2d�bAI$մ�q��a0l���%n"�.�n.�#;���>r#��>H;�3�_�繘Z�=�9^88��L�����ܳ��yĬ�q<�M��m�铣1�;)�$:�����#�����)�J#�����0u�2ǒB���n�RT@��AJ/�W�d�
P^���E3!V��EG��#ɼP
L�󲴁��R`�d(;B���`�5�q�6绦L�X���� s-�4"��S���s^$H��E�L�%�4Y��$��1"��><h��V��]"V8UI�ߞ��ӈ�����QX)'���ˈs�m��y��`a �8��)�.�-ͅ���8&��7W,D;���r9̢�c���oNj�T�`���Ԁ�i���N"Pc��G�~��N�H�o\�Z����s
ޱg�63���kVC�лƝey1:�X�n�&Hyft������^���~ڂ?���S%���dC'��f|����a�`���s_AHk}��8�L�����Aŏ��¬�L�I�3;F%9����{���H����@o>�P����|��Ӷs��8����DTA{�c�w�ѓ,W�
C�6�i]-u�=�����yQ�Z���6B�[� vş��AJ9�v!���c,���(���2UһUz�ք��L�zs�`����\0���&��\��NFnZ���'^Ri�(H�v��s����F@;�\�c�5"�Ӵ�t�vA�Q>=�J[�OB��jl^��0n��e���=0�q�b�>��C+t�`��D�B�,f��p�������i_��hn�����X�&��ǺM�aw����Ie$!���k����t(���L�d��d¶�\�k�)�F8�v/�u�e�S�~�P��R�O�"A��jLr�*"&�����6��B� �Y��&Ϧ#����}l�4u���U?P����
�`c��9�|��gm�ɻ��>�������{�}C�Z�_Z���������_ ಬS@(� j�Ⱥ.�����1K`O�g�� �����@�SP����2���\t����`2� � �b���J���q�������ˑz����_�I;_S�׆��B�p�i�L[(0�|A��O3�5���9D����Iș;3�.����a�ZCqTW��+Ǽ�����ٓ���\�=����Q��֝+/�= ����{⢭��y���bWH�0�%9����"�e�]k���J(��A�dQ�ګ��]�X[�\(�IYKw��B_���@���E��{�n���D��%�{T"��A�O;c����Ɂ�ƕ�gB�����8+�ՄG���a^��4�w}��P�)R떙ZVG �D��Pr��[Dh�y5Z`���j8��\�W>aߵ�T{���q�f3���D1���pR��@(g����FC8����@@9�_�����uS�E�4�}U���r�C��&�H���2M��!#�<��TiޡCp�¤˦Ei��& "�WXm��c�q��]{��̿��.�@��U�,~���"��)�!v��e��<�jl���qfൈQF���@?M���0Z��po���I�p|P�3Dջe��=�Ҋ�,>r���ه��8�6�U��eqyAs������=Rǂw�/s�g8�?
�wU�7��M�k���1R���l_����������3:���U߽&��5 X��+�K2&�����)*T�l�9�E���ev���5W��Ƴ�	��f���!�Zu�جi ��W�Lu����Od�`ۇāqa�&Ri���!8��bҮ�=��8<Hr�i���>�B_iy#\'*Y���b�8�n��p��T�\��,dPR�ki�&��Z"�so:�UG��Vg�,�yЏ�J�NJ0ށ�l|rBJ�̐B�gq���?@�}�]t�}L|��z#`^:�&�:��!>pC	P���-��=h�f�����)�~�3�N����sX�ؖ��`��;�6bo�$��&B�l��~��ƔI@Z^�\]��׎�K(�kG�c�'���D(�Ҁ����"�.���Lɟ�w#��a�f��ϻe��ϯ����YX� ������3��^�x�/�]))�A�}t��ԤnϖJ0��9v�O|��Փ�u�bt��r����ْ���U�Ѡ���ֽ#D�T��?\�[g|,q��_k�R�����e�)�Qޞ�].)��P����?u.��-�v[��g��UFֳ�u撖��bS3W?�Q�<��"0D������	?��C�����{)g�)���<)a���:0>K��9[ �!�`x�D�b>$�3�铮���n�e��p\��n�=��uIÂU'���ɇ��_����\E��ۃ�ٷP����cH:���'�47-�mJ�7ݵ��&���~�j�'1�I����,.����$c�q��B������:o3jɷ�aX3}δ����Ύ5om�٫����]���W�d5�c�@�EF��(>�E�ʬ�lF�gGa��d�������Q�"�>qײ�\�x?myk�\��ZE�xL�~�`	(y\9��(�]���x(�?�a�/�������k�<�f�>f����GZ#�f�
h�?9X�j���ӽ�{�9V}�y�!��G�����{Yܜ	@��ߑ�s��ގ�V�C�b��@���R�o�fc}B�bk"w���2��^q��{Hh�"WQ�yjÏ�����
�!n瓎���(�Ok�d{g�fπ�����A4�`߫�j�⹔m/��M�o��ĭ�*0�q��\�"x��$)@,�ѯ�k����턬y��~��_��1��\8�WF�1����A�?�Icf_�'0�h����^���L��2!a��R��\�cw>�������8� �K�j÷p����$+UccF�M������ןĒ�%o!�_G���㜬p1���/j3Q�����݀W���3'鞚�"l��6R�Uo�	r�j���~�����o�����=0�񘵗M'������}�����c1�J�Vڬ�A�s�v��xP�v��Ċ�{�������G��Hc��s��*w��C�>x��
86��W@)��i��ϳY��1=���L -��ؠ��W9E������!�M@O���9��1��%fF�~;��~x���h��h戋U�t�	���mMdE���v�OO��-M���e��_(رu�D��ɄS����tá򘱕�/�K����9+�Y�����Jm�=�vh�;� �޸����D��i~�6��� �`R�Xč�6Bt�d|2 ��������	ߐz
���gS�,��m�?����"�]�	:	��������텋��d8�F�7�Ѱ���m�>=�ƖQ�H��?����m#�ڬ��b}h�b̌(צ����bo��{<y7�������As�Ϝ9n��G�X���ҋ��?���l����X6ؽb�96=:�9z�yO����l���ޢkz�k�)ө� ].ů}y1�@�<A��DF�ѵ{Q3+�ӛ�3��X�/}^F�2[ϱy��ps��fW�6vs�9X�MA�@��|�3��f
���O���4L�h�8|���/�@����\4)�%*��&=x��~���;���kIT~�*QK0\�D:tU�{��*b?{V�|�d�V�EI�����C�It%ȧ��N� F�����X3^��Y<a]�^�}3�ŉ?�S��#�S�8���V:1�H@$�"��7D��7r]�bQ/9)���D��yNB0[F 6��WY3����\H��?e�nި����Z�}-�m�ۍ�<s�0�JkaXx� 6�Q�¶�`i4H� 7�,oπ���>z9.9�+f�u5���ʀ���E.�OpC�j
,=�@u�tQ�[����!D�&*�6�!/��A�{�wy���*���}S\�R�x(x�]$�X��
��.!���gzd.�v��ޱb�z�������h�5�?_|V��v�RH&ޱ��k�qWT�ib���S����0
t�<���F~ng���	h��I$ԫ�<p�:�Eŗ��� �u]j	ڃ�3Am����\�.򼗔}��Z>���_ۆ�BB��[׾�	M���&��B�� 9K�pz����E��,��`��m0���U9��I4����|iRP�,o R���W�5�@���M�
���'9�qW����� ^�Z���ԳC5��q�Q骧��s��y��Ñ��d��&B�'p�0�p�w(:i�`4gy��_�+Z�E��E���6�I?��l^ɱ?��0��>â�,"��a��	��ec�v��%�pDe��d2���:9{݈��f�7�!�@�B�� JT�'��4�{��n� �IP&[W��E�Aһҫ�6��UN�غ�G �+�g�c	v�3E��B~T�ݠA��z�$��փ-->��Kl�`�]-	�0��=�L�^0`�sEv�vHSŽ�0����' ��\K�M��.�;!&��EZ��~ҡe��۸�1�U+��r����9�iP)A�`N�	�3�J�����nV��1fI�|'w��jڛ�c����H���W	�F{�Hl��_d7ja�0Q��5[��]旆˶өH[�$�_d��
z{�~������ԄE���=�J"o�ڂ3�/ xR���
z��'�ݞ���,����?QL ��/��p�@��ڴ��z����5~.l�E������p�J�����N�0�m�	yu�/��E�����j�t�������c);}l}�¾�������uO�b�?�Xt-���-4�sh�:?W�'9P.���CU�bC�t`�CC6 �)e�T�r���U�!�bW��ɑp+F��k���]�R�oe�v�>e�jPٰF�6�6�_¼��,��y��vH�����dO��(�>�ʬ�l[6����-�ג�	)`@9L�������F�a�J\e��y�C{�Oh2#�c5�W�Y)�H/LF�h���D�~'^��^RD&A��ˍ��4)Bǔk�b }~�G�������93��m
�{��S8~���/���$����w��(�t�pU6��<u���ᙀnW̦_�b�F2~��}Q� 2sʂ{�q�X�Q=�����-f�z1�A��#�B3��شz�A�>82_B���J_�|���F9U����U�{�P���&L1�h�E?���.�OK,Va �����㧮rW��}vi\�-8����6
����g ���[ =������{2`{��㛱]�n�IB��W�����4����=o	�����+	{X�D�S� �!s��b���T~�LF+Ӥ�5:�`�iO,�=:��oDaE��>��1�u��`��/̶��㚣�č�.E8�|B��!��3J���T�t��K*��(�����)�w�e2�}7����9�7W�Gޢ�:��s�MayL�g�!P���fԣZ�*]���ݬ�4�:�]72�wV5iī9�p-�/��&� ��J��*Q
���w�f4��/��/A����̖PTa���&վ���-M�v�՞_# MR?f�D�0!l��h$}� �WU]fZˣ��&�
�����ĝ�SQ�<�C%�L�u;��3�`ߞme�/��:�4SHQ�m�#I��=�ޑ�5zIw�������u�$��i���B_}���,R�hҥ-{ 6^�}l�,��I0gH��Ne�k/�1��Bj�[���f�Q��L���=D#�z���m�nrf|G�*?��*�oB����A�A��8��ϧ�|�ї�~"��j(p��J��U��tͮ�T���5��)��ʅ\���S@�p �O|.�8�4Y@�����������7�����F��~
�!�M���D��_��7���ʊ�:G�&1�s���9���w���'��w���LN�T0D9��S���`��V3]k�D�o�O0��ୀɰ*͝�	�P��ȋh{��ЀF����
's]���.-!���* Ȓ#�o���̝��0Wᣴ�Li�:��?�F�~5Q��VyB�������	r���7ʒ��
$�MV~O�� [��Dp�q��/�,`tF\�2�g�p L&:8ѿ6��FT4��р��m-S9�h����]�Cx	&�Y��1>�J�E�Շ��!������0.��{������aT2�s��v��A[�8��W)t@J�Jx�� "�kX��"�mpGU�y�.%��*(�Se�Mao�7Of�t4^���x�	gz��c�����XCn�J@,�e[7�˾G���ɰ9�2���� �h�$�dqq��9�x�LM��rI�p��k����Lܑ�	0�K^T�$�H�+��IX�����y�T
����Y5W@�WR���`�����rIH�p��k(�O�4��.�ԗ[��1��d(����'���ѐ�a��5_m���Q0��NCk!$�����Crc5�J���'[6
g�R3eO����t�'e��-x��X`G�"���P��	p�S>���bnK닋�r��a�b�����'��!�Bf��<���HN��{d@�Ϯ�¸R�a����u�� );�A%�;W�>����f}+�l9�9R�ZU"���F��>�~)��Vv�&m�݅��+��~��=w���]Ҷ�$�E��˻���Y�ˤ���irϴ����Q����S��؅e��.����}�Q�l>��lqO�$^���33�w F�Γz��)"�RY�h����Q����ѐ\��Q��������6 m���j�L���G��� H��E�5IL���zѭP�T�  `F�A��I7X�
�LR���h�h�es�?e{��ٛl�jf��Ȩ��[;��Q��92�3�sN���2�&m��H�#5�]�=}�'�::���n����LC=C�C�>}���7��|���)P�����t���dR`5⎿�eDm/�}���!Z8]�B���҂Jړ���Qj�B�?B'x�<��bs��h�tU�t��A�[�Vs���4��ŀpMy+�t��(Tß���d�:�O䁁��'"�<ч�U2~��^!Z�u�3�r��x��o�( ��x�{Th� �!IWQ����@H���]PȒ�9�z_{��%���q3��uK����ߪ�5�q���U�aϝ��SB|�c.e��~�u�_0��O�0�I�$�\��QU%G�-�҅A3~E���=R�2��������JZ[\��]�C�g�R��B������G:�����ًSt��[g�7;��Aѡ��WkZ��z�ۏP�wtM��y%u�/�!*�X0X�l���HG�5 G��+�?����#{�l�7(���j��ym�<�;ߣ�E}���^Ta���a��b�w�}pEq75���q�~i�جy�u�:z7��{Y�G�������(u?入}�4�ͻ=��U���"��n�i{|�**�o~��҂�j�vz|S_{L�����Q�zx���y�hd�������0Y�x���S�|+��
?ʼ��.Oƽ�D�1��o�}��N�A��Ԙ���;x�%#��������XKKK� �>�
�%�+]�������]�T!�����O��9�!�+Ƨ������Y)���)gʆ(Z"6���8e.+a�^Y��$�k��ۋ�ҕ�u��#]_�8g�K��	��Q
��U(���	��3PUc��o��'q�wd�{Μ�z���V��t"?���[����vYL�O� d �ܮ���L1
!��$t���&��[���K��[H�sJ4B蟚��'�V�-Ф\�x����7��ŋM��0�;}c1�\PJ�Me�\j��4�f(n�Չ�n�t/b\�+$"��*�|��w�fI~%�6��p1����bԵ5���fr���)�3�r�B�֍���3��F�2r_�V�ɬ��|B��K3�1�	���%���n�]�)�w!p�\;h�ԑ��Vv ˜�4ۇ���'�p������f%�� .��U��R?p��mĵ��i�����o+?@>H��Ey��4�k	W�w	*�9,A*����D]|���_���I��(�Z���g�+�D��X������M�����05.0�B$��F�Zl���!�"�� �pOC�v'���#� b�Nɏč�C��V�"�S��<��;/N�ҟWi�`O��&2���vsu��..��D�}2_���=�2�T��R:��	y{�p���Vg9y�9�*���.7�a%Fb2��L������~�yO�Z�<�$l��/OA�M�v�7���0�ne����D@2bߴC��$(a��sİ�KS���ȉ��Mc���̾i��vp	M�{�$�k$v�H<~�j������c�m�iOIc\A �(>L{��RW�,,��Vq��M�Ud�FY���B@�j@���w�|���,dd���Ho���r�4
��X�x�?�R|ڵ���U���-/���w��Fx#mf!eP�"�@>��z�I�b�]1��Q*@�$�-�+G-e0�����у�K��y}�ߠ�k:e�������dR��+��P	��l���<�Щ�<���Iw�N�2��}�-��.���\��T$LB,��5���+�=}Kօv2�|v�M�Fʸ&of1ٖv�X�p��.��	�q�-mA�/*I�[���gw?�wk���Q,;�u8�͚7]R��Y�1�K�#uw����X[7���@P��`�2C�;�7��u�y0� ��|�f�D�����T�fZ�u�����b8�Wć�M.��5��'wR�-�	ԮXJ��֝Y���J��&mqt#C���a��wp>$d�/�̟��XD�{N�3��9���W6�|cZ!���8�b��M�	��х�y�WU��]|����5İ�^;r2�l�I�X�c7E�y��~5�ϣ�*�i���`a���6������ھ���A�=��*�ܼ��wq����yf�;	��.�K�6q��t�s��8$��eqȚ[!:QRx00z������R%�k�<��E�-�9�Q�X)J���j�DO DZ�i�?�%˙��*����u�8\#S/�OQX5�R5�x@�g��M��$��g`���
�N@���2z>{���u����@MZĂ�cb�!|�C�%�(�7V��A$�R������/av\�^n� �����l�����AL�z�D�C��ݬTN\y��@=�J��#Y���rtG1�;tO�E�m[����!�Q96��~�ǜ���'�1#�pb�-t� e�0֎��fN�k�K��� Z���;]$�q���1��.�M����`��Y��S�'�ӻ6�+���m��r�E����gK��r� �k㒢��b�
�̈�Q�"+��m�t�y"�I�I����n��r}�rH,�/u�o��Rd+fP@�B�R����+1Rq'�񎙹�WOu�KՋ���&K���^[ϧ�D�Z��%���
�q�y&�ϊm�t��12>PZ�eH�c$�����$p���]A��o���ئ~8��H+O�&A�J%�߻T����M3�^���x��]Y�����AK*��7 �E`QGz�w�������ͩ  W��i��2y�qܦ�Z��uF(�(��^|�q���� ��#�=��� YC��%�r
��^������W��9q�A�w��L�9O��"e�mO���S���?�
w������`ܢ�� �MD��H��r�v+I�+"��]���g��?U�ɝ{���B��]4���K�0��	�Ys�%ѯ�w��q��Sp��a�����/�Xbw[\ |�h��HT&NL��	),��t
����T���" �HKwva�&yl��+�vf*-���1��|*�5�UX��+��,FvaVS{������_��1�c���ªˇ��$-ww=5��)Nv�M�Vn�uhک��^6Ւ�>I�'ڠ�ϫ_RY:4�KI9����:+C�TO雕Hi˨l����>�4�7# ��ep񍗀������fĊr��EWy�'�������-���
����q�}�P9#OJ�Eߗ^o���y�{����"� ��//�38n�ˋ��T�iZ�b�
��"69<M��ނ�>�F�nS����J��5-m7@�����t��m�EI#
�H_����A}Q6,�����3�����N���0Yd��cc�H�^���*�B�[�����k��h�ھ#@��.�=��p�Gjs={�}�M^��c�z�/��\fo�)�'�ꛫ����M+��As���~V�Q׽�x۱߭�	�	�~m/�9�m�!�\���l�1���I��Bފ���L��0��M���-a_���,����7)�W����ݟ�E?����JH0V@:{�chd9g����(U�f�K"�2X�U}Q�q�'w釾@�vVБ�5��8r�[��8i�q�ş��l�sCT��t���Z?(�0j>t���ZA��տ3���\�X�r#~�C�2�盙�>����N^Y��m=6]�@Yw�2'��]�� o=
�^�����is�%'��8q�SvB��cA/ө0E�@�^	{K�_^��`�X0l�\Y�R��{�m����������6��7u�p��/�����mg��=�Tt��c�r���ď2g���Mذ~_f��QE�37P`��4D��s��Ø�օ�h2�<=����< vV)����_\���q�"�~?�#�eN`��K��j�j�9����"2v�!�hc�0��7-�X�4]a!7�z�/Ƙe`	j����=��B�%)��J�0Fj�D�xq5�V�� -8��)�Q	�$y/���b�Ȍ݆��Č�mr��0h��3�G&��o�gsg8zJ��>r�.�]���*����P�"I�ʵ6��j��ҥ./T�96]�ф'Xd�8���
ɋ��l&�eҨ��G��L�A����FF/\P���>p
��&��K���Ð�qG�����}qh%�
}�7�@d�
8�e�'ϖ㮥�{�j�	����C�FK��G�J����?Y�����p����\�x�8K��(�5�G+�)�qh�R$y9-��l"�0���������i�#����K��e 9Z^洖z��Tl���y�)�ru-��2��C��+4Z������W�lpƬ8=��G!�zO�-9�s�[:�bg�@7^��������x�i�ݕ\��Zxe?(b��6:L�ŬZn�G#D-��*�>hY8ܨp<�34��6�w�+��hj}�e/�ѻ���A��ź�����
A �,�l2.Z�����W�R.��%1(ď���j���ֹe%w�Q���&��ds��DS͒S�w�Ő�A,7��w`"��^������`��%���>��u�
c�L� ��Y�1<�K_9���#�u�}<op�PS��Y[m�o�K���ҘJJ�ĐX7 b�_�c�n�ˁ%�%���|�#�� _6�?T��-�ɜ�Z\��T�)��c�N�q+lNi^�TUܓ'�l���gs�_����͐Jt���>������T��]�E����h5N���PS�A?�CIXN���}����SBȚ�a��3ہ��&�����)~�%&�[��x����2�O��=?���<L�џ�j�JR�`M��
�,_�b92P�l��x��y��.���T3�N0pV�dV>%�M�L���-����-��<Ӹ�"����Cv�����s����3!�<���X�ثR8�:N�Z��&� ��ۡ��X���-)��0B'۝��0�I_�n�m��P=��u�"�W�w�����v~8KK��5��qJ��a���Jẻ��~���(oLAh��{�z����q�{E��}��PFR.i^up�ƎaGz����E~�}�"/	��ka����hD��k1(��hQ>���4����,tf�x�����sV��}wlGM	0�0�L(��J���l�c����`U�]�d�F�5�n��#�M�Dv%hn����U$�8���
kT6Д^Pw��d��t�p�ʬ`��c`�ncE:��Z*N!C�У~%W��(��`�`�N:�7[V"H�Q�2�L7�!�J*"Bm����by)���j�#Lx`� �0���|��9r�c��0h}¶�&X������<=`pTW,�g ^�wAU�bf�Cf������}�=Iy\;=������G7ڌ����tX*�x��Ѿ�Z���<ٴs���I޹h�m/��I�f'X���_�S�]$������|��<xJ�\T��W��uбt�$j��r���П�i���ɒfz�'\Gth5I 4�C�_��^x\
9z4I�+B����O��.X|3�>��d�:���_�pQ�����N�(?�-H�-��Ix�m����0�������w^����l�����t6�q���^�o��R/��mS�����H��sY�ؼ#��ǈ�����*�X���Kg��C=W9��������b�5�f}>��9���d���9�N�	(�w���Ϭ�]
�Z����������iwR��d��F��̣�+XEϙS��DVj�o�;��f�2�*~�ᆷpJZ��Q6gI�-0���x~�;��~�fU�� Gq�\Jˡ�x������Dw�.z8_�o6/��Y�n�Yko���(ꊼ~�7Q���#c9��5K7g�Ʃ�U��э��;���US�^Z����qo�N� ����Ӵ�[&�XI:�s�(N8X���{y��V�P�t{Gns�,�܍�Cr�#_Z�hg�IKDQ ��qݏ�=�NW؆��ԧ���Th�򒿖ҋ��F�ڛ���Nl*8C�����t��1�-<UN
"�/�����J�'�R|�2��]�>ق���˟���{I��u�0$O��Y;�i����8��M��&�.G+~K���^�;�	��}�C��4dn�Pv�B3x�0��1x''{+n��I*:&~�K�i��	~��4�xܕ�[��F�hH(��׷�@s��S�g�.�=)��6_�`|��@$��؏s�%�k�!��orUGa�yNh6��{?]b~}U>���mߜ=����K�M�fl8��XZt���d ��7&�
�d��!��z8HY�j����l�D��G��xؖ�
�+7�M��:�*%�3UQ���{Q%�Iuh��ٲiTw���2$��E�3-�E���ݝ���{���ڏ:�gh)>W>��"H{���}��h
=ֆ�G~�!}�>����{��T��WFa�X1���m�]
?J�g����@�s��F�bWX�!r#8%�������Ҙ���CA?�hPY��*���-���@�2k���E\O~p�-���z[��k��] ���N���������X�c�D]�}#�D�rd� ���y�o]��Wo˸[�pj��m��8������5��x&+��KR���/�:� ����3�G�n���%9-��9�Ϟ�Y,XeH�U�e�rH�Y�ښ���>nzb��P�8�϶#U����-MAv���״4�?�ɼ��^h�Q�po��|pX]�C�0��CV�|�Qɬ���?h��;��k��=|�&Y"���}�}S�R9�L�9�Ez�T��%v�x��i�#>>��Ʌ~��!0�Y������e�+�5Y��h�u�cuԒ��񖓱��{9��dͱ�#x�'��i��_t�8V�>Bϋ�7��]�2&~�=X)�8c:����u���V�T8���J��}L��b!pnr���o7~c�?��?�C��Ԥ���,u~�c��Dl�Qj�m�ʋ6/��$`E�Ȉ��o�^���5I�O\J�!,N��@��d�	��;���c�i�8\Lx��~^��L/4CZ���d��P¹y5�l}-�Ш;��NB�w��e9nTZd:�6��"��) ��GG�6qI>�k�M�N�@������pe�k�i���	�4��2t~O]D'�ψSŋ�<+��1l~��o�r|"���g�o��F��@��G$Ǥﶼ�l���p]�B�4iN�[𗘾Kj�-P�/^�O�?�����=��H��_�ʉ�2��յYɃ���"���o�o��	��u3���� /�Wy޸�P���</Iw�S�
:�5�|e��`<0���X�ڝt���n|��d%m�P�����3����w9���ʅt:�x�aUI�ֱ��o��>+��*I*�8]��炬?��U��!�ۗj�`Hn���ע�x��B���7��k�\��w���<yD�u-��]~%�Rɀ�T+Qf&��Z#���3�N�l�cSo�D�y0�L�L��cA�6������hٯ�a������B�V�r(K��=xp��U��>G`��Yfٱ��&�m�y��N'�#����V���k�n���a� B��,�ңF�[���_|�wz�
r�zt����4���lIVN�����aؠ����y�a��nO�xB��GӨ�|���T����	�>7��G�p��l�ş�7B��<|w�c�h�6�7��ew�P=
7�~2Ȼ���i�<}Z�6Ϳ9�5+�f�1S�UFCZZ��!s�H�j�����b6��&�s�pz����t���5A�m�=da�!m�e��z�^��?o.��4�W���x�tt4	��U$ov$O��oD|���7�������R��1�2oA{��R����"Y��X��x>
������+Ã T�_�!f�.O���VT���A9�}w$�Zk�,�+3��	9V�E�W��.���m��m�*p�r9�T{|/Q��*�!�d��_y��c�+w�N֝]����a
�i6|U���P]ȿ��s�7r�Z����@��Ooڍ�5������~=+����54+�Ű�Vѧ_	O-!xy�[�f�=�i7t7��d�%"��&��C�yO�?^�@�ּ�)��9�2�ɨy�mw] �{�%���c~1�r3�f��d��[�FO���w��Z�52�����{I�^)�] MB�Z|UE)�U���#��)��s}�|���u�9F�$�X�R�˿� �7�x	w8v�<���\�G;�-�Ò�ow����ʎ�}]��7�眴]f�Uc�<�f����0�8����H-�M�8ò<��VK���m�
�|����
2W]�<&�) ���ޫ1GG��#�o�b��\���ŧq��P:�&8١�6V����q@��1���>���`Srk=tN�l[�8������j=�+��b��W2+_�AtG�[���w���!ݬX��~l׈�G¡�&��ֽ��<�Y+�^�8�0�r(8L��|OP�I�Cy�JC0���R<v6��緞yKE�+�h!���L��R`���<�d�����|��t�>� p���DU��%�W�`��M.&aU�7����M&�����1�g$�7�
���:`�mo&�g�%.m)��"�{�-�&5�[I���%?x����`t�L�g6��:��bG���������yΜ�,<W��H�<R���J�\^١6��9-����+
�f&�{�,�*˓�|�)�>x� ��Q��XX?³M>��|Ҽ?Y+�@Ѐ�H�O>�s*�M��Ԍ^���*(��S�7���ȥ��vK�����4�O��c_���b�*�˷��͂{�%4P�^c��DT����?D���#�����l$s��7�� l��3SnD|eQ�R^"���#�m�)t��_��ss���h"Nœ�����e�����纳� ,q�H,:�ܦO�M�<����y,�g驂���f� ��7"'OOC]w����Rj�..�6��U\=6�s���)hw&k��������+ꩴ'�S6�?"OW�c�,��2z��E��򪦚c����X�:�A^6�#���~��Ĕ�TufU�WƖ��CN�,���O�U�m�#A�i�(����Ow��1����P�q*�����t�z�|_X�2">�-����y�$�\5W�_1%rJgu�_��,HkW|J��o։-�K�l(����[=?��|_ơ�k$�OI�Qa�[�Tsp��!��ͽ$dIg%�B
U���o8!���o� �ϊٝ�J�꣑�2aL�`�~h����N�H��8�4�ա�%�~�SO����P��[A<2���?i�zĺX8
0��W*���a�����$]::�EY�\�[������W�%4�(�#|V�bS��Ӕ��
� Jц��z�����Q�^��*��� PK!��ޭ���OH������:���u�H%��M�M�aWt#`��������
Ç�#�y����*\�G��Ak��UG-�1�M�=A1s�Q*�g��	`r����ܩ��e<15�@3�/��KX��@f�ު�ԸH�t�_P��{�t�b�
�a�{��l�E��!f�N�}4
�t�=����z�1I�q������O��c�)�IЍc���|d����NuYc�?����z�����T������Iݿ�K��8t��j��+n��(���k�8�N�N�Ft/2�l��ٜ�R�6����}	�iAР�+��vE#?Z����{i��ɕ�, ڶ�U�FV�z
��SY��CG_n[�3��fP2;��j��6Y��	�����D"O�������*dY�=fc���`����
k����d��Vmx�t�(B�V��l��9�Q_��#�����H��_��E7���@х��	uݶ�<5d�wxi��1���r���wm҅��.̕���q�EWc�U�hk		��7 ʔ�-���p@�P^�0͈���1԰i�!�aN��ĥ޿�ҁ�`�W���n��uE�G�켔K4���?רgyIe�h�Tuu��\I��{�Ǫ��b�C����"��\0�|���R�[-���\ynwc�Hr�̰��h��l��2Pz�3�y�����A�<��},��(�N����:i8ر����03�����? j���,�w�ݣV���n�)96[���p쎄��#b�����G�q��T��"|��׹��PiV^�l�_t#���ŗ�[#?9�-���!��͡�&�~�������QR�g�%Th��ۛi_�%�B�l�v?��vp%����%��"kE��Ir"�_���aM/=~[%k�v8g֯`(�#|�+�!(�v�0���zV����N��;%�k���9�wXL+ �����l�P6y�T����qP�&b}�hy��5�9T�`��
5���ƫ���Q���׫�B�L��G���L�2r���k�Q-���z��V*�'1h�'P�S�Y�	+ �5T�{@�"7.eϧ#׎8�,6�=���ƗfH�9����}��H�1sO�I�3�]�R��x�u�_8ʫ<F����	(�Y�����B�U$[�F�re�w[�����N�g�tGt��s��߾F�%��\��}I��Oֺ�@L�aL�R�X������.vm�|����O�>���
憰�n,�.��:L��X~�o�﨤D��z�M�������}��v�]�;u�_�$����}�#vШ&$17�?��m�ڿ�k	�b�b��@�3A���Ӽ��L��ՙU(��/����'���a�z���5%��htk���Y��HN��	��ܠϜ�� �1��?a���7�n$]�
l(�����6�IxW�08R���3��r+�?
���60bF���0�� ���e.mB�O�č���*P�%��W��l&��3�L�v�
Hgg���6�p��ⷉ�vz��Y��r�	�1�<�sb���W~D��k�Q�e��@V�=�e��	%��a>v�g˪�]3��/�LA?�	`n~�7�S� ��q��-o�5�dj���/ߪ�S�O�è�~�O�m�]�8a���sv�h�3��c��%�[3gk�v�i<N넭���z����̥84�EJZ���z�Y�.5�1+�ْ��ŝ��a��|����D� b�.�=P֜v��+~�B�\+~�1�T�M&R��T����㉩ ^��b�&���.�tr
�%�Щ��k�E�v S�R���`���T7j�/	���jƩ��4ql��G��9I�R�]��"2+#%�l����	��8[��:9���G�����*/>�`��T�U�7e�plG]��@�b���M�l�MH\���0��ZZ�����3���jŎ��x+!��b���߄��4ղݑs&�o���GZ	I���"����1��y���3�bR5�i��,O�D_ܵ����	�z���+��u4��{���Z	�d����\�+o�4oGNg$�ӯ�nי�Ùv9�N��[W��n厽�l����U��f�y�ˍ�ӻ[�eAP/��װ�9�pA�Q�[��,�NB�bw��t�l�,|�c�b�̡�q�0e�lt�l8-Yd���%1a)��@��d崀ۤȬѢ6��~�AH�ţu���t�G���N0L�|���g2D�Y7sa����c��'f�5��ɥ�n�b<��SQ���p�B�slne������3pD��3�l���f�uZmH������O�~�&�"�� ��=�o0۬�r/c�4Iݾ� %ͱ�^|�P�68�L�JJ��Km�r'��x��e�2!�[]~��3����eR��qJ����t��D�1;�<�<VI��G�H�b���O����Ԣ��0i�'|A��3�A���M'�A��
���N�$�0BYx�%@�W2���F����=�~G��d��`�u��s�Ԡy�Ѧ.��};�_iٟ(_1,��yҎ��L�ǯ�A:'4`{Pv1Tt2����֎k����ܰ�;�@Ğ�%O�߉�o�rc�*k��K���JM/n*�M|�l[��3u�)����3]���Tlƒo�Cpߠx����ox�� �TQ�>�}kd
_����f�b��T�yLC���N�^��S]N�u	p\�=�G	zk�<���)����ڊ{"���։�*������A+��q����Y������`�
N��2�啱�2�3��o���E�%���B�DÞ�����-|3*��Zs�^J�
�rk���	W��Դ&v�l`��@�f�?�e�;�*W��$�P�TB���F6�h��q�M�?��e�I#F�͕�t��,��<	�(��(�������f���'�8!(\Z��I�s�s\���ΦL@�LLxdIrcI^��(P}�;f������ȅs�������n'����qL�g�>�a��1n�_i���pq&&���W[���ׅ��m	ےy$odu�FY�N\���{���)@�i89>�.�]��^�%L����FD�W9������\0J�ش�P0ؑ��+ZN;h譆	�Pqs�[���=`�R�}BR�'��h7*�:�M&�gC�٠�zw�i^�σ�y���}��ٶl���%��ٳ �
w��%Dm�BjTόu��<jhj:���������ƴE�y?Ux9�b�̇�X��]��L,1��
p� �#Ĥ?���4�A.���M 1a]����*_�oV�5��W��ь +"�����aWDBY�����y���\�ժ!_R����@����`3�lѐw�f�����T�&��^o�����@K?�f�86�Ӭ ���WO����Q�l(�U
��X�a'���U������{����Aq�	oӥ�G�%)���G{��^ԡ�+]o 
�W�ah)��~eW;i���
c�{0���~JTnS��EA�(��m�Fѷ��?g=��.t�"�\K@�%��}���Ve2Kژ&��-n3�;Q�q-4nq��l����*6_�~ɱ͸��bnb�_�;/�:c�5a1%6���4ޯ2]6�&6�JTHs�@qo�*�?/MI�p�}��X������� �K%ʥcͥDN��0.��ǖ�oKG@a�fX@��`Ӗ�U�}63v�
k�' ��	��,a�䷇��c�G1��Q �Q�.��g7���D�P����X����#���?��?a�{}�s.M�ī��}	��ɿ>?��5��:pj�bRD�ݶ�`��Gxq`��JV7�)�k�W�L����c��K�{$J�&�(��H%�=�B�5J�Log��S�ۃ�퇨Z&S�����/��=����J�_��yw�ru�)k�^���"�S7��� Sꏰ
����n���k�F+|.��e�r1��lQ�#��Ԋn�5*�*������̝����� �µ���:�bvHRFWɪ�V% �����`|)�*=��+%KI����w�#wM
w�����D�,�e�7r�_�Q���ސ��4��ɵP���ǫ��y(���˰x�RsT�����>���O ����B�{�o�!�O~�
�fʒ??"��*q�8F�q)�ȟ�X��I��+�����N ��q�?���w���n���6��X��g 7n���)o�?v1������o�}G�P4��yWgɧ���$^bYx�Z�4��yF������՟3��2��YȾ��&� 7kT����U	Lx�y�t�����Fh͚�����(�lf\.r[>���"��"�c�P��`��T$��Ý:�S��'����}J`����o�S����pJ/�e��`�QFEV|���<�~�_	u�1q��r{�0I�	�!�� ����/��4�]YG m��g(Xh��������W�/I�����|Ks�[��[��]īU9��^����x)�����B�
����qNg�/�'�fxE߁�����`�ʟ�wo�n�jc��8un'��C(�hX�{�<	�s����ΰ'���h��`�ʝ�?J�9W��z.f��\�_���(t�Sra4m�1|�7re���.�x�����^�����j0R.ӌW���|w��\���<"�%N��qcJ��S����3����{���+_���H��,a�}3Q\�I��0K4g��S/�o, �0|{�ؤ��6v4��U�l�uJ�Fb 5f�|�K�&��]ղ��'�3/py
�Y��!��vpR�ͨC{��K�؉-�"Li׳�r^^X��#�}L��h!/�B���>Ԧ���#`-d�=dV��k��:<b����~� ��I�K�!"z|>h�ad�4�^��}�<�]�7#�)��H������W�sd�=m�Ρm�z.����-�0�P\�(�1ȧ>|/w���4�2�����<��H�7?��7��w�Y|����d�ض��/8$�u+�f(%\yy~: �gA�%�8L`8ք����k��ҿ%!R|:����K��4+b"��x����H�|7]�A!KqP;�ug�oG���Ό�Ƴ���Y���(��0��@��-v[��2��mO�J.��"-I�9��u��=ܶ�%�P��=����.[e��#N}J�
�A%e� �n[\�;O^�e��+�h䫖h�'�o@�?5�%b�"�3���<n���6��a���<f;F�@w9����Y���q����h����I��䡰�8�x{e��ϱ�̥�0�.�h��Op���h���6�#Kz���B
�����5y���e�^F�{���Q��[���賁�J��vE���9G#ij\��4�#~�2�3��kb]V�W��I�=��E�����e��}�\b#��h^��zdӽ�	xhyըY������/W'U�wy5M�ȶ�;'��:%���P���N���N�sk|��n��\��&׷7���v�L�l��&��ǩ�S�8���#Q�c���6�h3�A��O����B<�T�|��,<�"���R����D�`��H�;�)�{u=�K�*$x��� ?��O|�JZ&�#)	3��'��r���X �k�$*��6���e�E���J��+��a�֭P|��묗��S��/&a4go\�U����ƿ}����N2�Z�nɋ�[�C�gbq"ޠ��!_4?����a����D����J�.	VL8V��h�2(�.�ud�a�rV�m�d��t��N�¡.#(/����h�A���U�&�9hk��l�Β�av�����,�ab�8%�j����*�� [2S��G�׎-A�Ap�M	��K�~�(��WQ��N��$��-{�1��a0T1���%�%ձ���6��9�J<�%�#���u�\�,�f5�#��d�9���x����5�ϓ��g�C�P�����1��EN\}�i� Q���b�.�Q�NXnA�cbc��Vs�`�� Z�}-}#�'R p#�Q��7��<�<'&��J�B*�U��׷/H�q����7��ٗ/�ZȕL���ĠRV5�}Q�c��w.P9l>�1��,�#��2�.�F�b��t`�����?����}5zp���6�>�>&�7c�,"�'�ZBM ���BQ���p�ܾ��*��a�E43�pq8Ϭ��"�����f>*e���yͰm(�����S5�-�u'����^ � ���킶�J�´�|=��@�������jTX��ċ�k��$GE����~U��ȳ����}�lL�R��d�L��r&o&���������a�=ؐ�޹9��야%v_���(*M	u̳%D��h��3�N��L��8{�ۋ�h��F���<R�T����w*F��w翭���� �L�b��;��a�N9�}^E:��B��fT�l����]ۘ.VU��Q�_����'?�n�\T�\�PX�kq~���ͳ���c�4�\��`�$6���V�o���#2����M�%�Q��W jyF~���S�VY_3��o��)85=� �}�?��c]K-�"���Ɓj�m2K8�u6��9uƾCt}��;j7�s�N�����`8���rS`�a���\v�'���"}��u	��;�]�=���Eu���ɰ�xRN��O4��/�?�4�R��4��ý��[-��;/M��~U���1���4`�S��j5�"/h_m�bu��7 ��q�Pz��e�`��-�!ï(�V���8n����C�l�����K3�e�Ɏojؾ�`�#���.d��01s�`PG ��;Tzcv�`UR��wd����)or���j~p�H�N��܄(�+�J�_�c�=����Vz�����)<iGu-�"�.����F0CZ�x����q�gN��w�r�V� ��K�J$��3��Yk`�L~ˢ���"�L��?%M��mB,RR�l7�AH����&�veb_�G���W�X��]C���g��|XrM�nJ�p�Vy(����*0
eT�������R���3~��DZ_!��.h�U�_���vk��Qk�� �6�O�29[�L�#�K�I�M=���o�v_���c��ߣ7�{�_�F8�
���������.�U�� v<�Q��C������v���×��p;�\�L띖cPG�u'�r��g��JOz-ԥ͞�鋼�N؀�4���(_'�S��/ϧ��\�2K<�WT�A�^m��OcE{�������R�	��![��*ks*-+�4eN�a?��zޞ�ą|5,�	Q"3v�]{��>� R:�|4_C�4rRx�y�n�s�Jc��Ѧ���1�;�c�=:�z�n���WX8�MbR*��R�>$���&k�':����5���#��.���z&:nA!4u���`�u�����pҠ�)P��&�[�WlZ���_�G}ʏ:�EGb�`B"�])�E�@�,&�Z��T7�p"�z'�yyNfok�̮�´�SX&��Ž�co���żf�h=G�F��6���z�Ր��A֗��!vO��d�����/��
�D����T.y|%����T����^�l�0d�9j@��%��$3�ֺn#X�}Ջ�%(�KKr�����>x���l��N�����ڞ���4��m���}�6K�ׅ�>T��_�����&�E�z�Q����=N:.���1/!��CΩG@���9��x^AՇ�ZT���I0��bb���p�))}V�
�5�tY2h���1�2S@�Dx~��S,u�7���qG��5���z�� �ͱ�����Ӈ3���c^��K�ܺ����Y.�E�m�}��ۥp�Z��M�i���MW	����>6k�^�?�KY�3��V �yWVs����v�CN.
h�t��&�k=����k�dv�8��C��e]�|K"�������_l��g��?��VmjsجtA��XG��;L
J2�����g�q�>`�G&v?�a�)ϭ� �x�w!^�����N��������z�uW���CWD��Z1+�0���j�MY�"�_��_غހA��Y�¶J]Vl╱�j��e�Ә�pJ]!7���t$WK�I�<H��Ԇx�;�fءKnf�%���Yk1�P���K��W�> �8��J�K+�G�_�S8*��4	?vR��y���n��HA�m���O4�b�g���3�J�r�s�ϕ_v�ms�l�^�x^lVl�a�nM�m�C�7\{�k�.m����l��in(�b��������j��Kb��%_������6�j�V&wnp����@��q�0�{37�8���"��٦Fh&��z���F��rtܼ��En��LX�R^K0OX�'^���}7x�,���[�=��Ոb7��
*tm:�=?�O��"SnN���L�q��U�Y~�_�h��S�%X����j��6w%�0���D�oe�����]/;
9Ϳ�����S���x�m1
�S�B�Vɰ��<D돴Qg{L��q�E:�V�ͷ��'Ψ���4��C�A�'_��Hm�M�	"%۰��^;���J)HΓ��8na#�E����g��:|�<�#iX�A�5tOqtkd��Ag�.w��G��>b���Qԏ����|�?�;L��j!�������e�P�oZ�����ݲ�B�w����t�}'�$�t���	�>3���)^R�#m���\o�Q�Ns_1t�����tEJ#�	���)��%N@o�� A�hv���|A����,�p���^/�N�ί������2��9�Bx?���V��\�_�w�2��1́ߖZ\�c{�9s��Ga�05LN�uqg�<X���ȍ-�H��>�\ƨ�����ˡ��!�u�%�/�ڽC�H������͟י͌�\+2�w�����"\�=�
o8W_ !�r���y���Cj���E�+���t�9�5�%������w��hY��v�9�01q���Ct�)@�,���h$��������س�M���y��8���G0���w�	�����T9Oi0��!Eu��vȹa�E��*�&�|�U��F��7jz}|x����O-��p9�� ���N��§�#%ȅ�"����-����h�	1ZS ו�ļ�?��c&���m�����D��Xj�t+�s��b�7�72�jD��TJJ��1}��H�����������A�ӎ�\myk���jA�#!Ң�Ih��0��N��H���נ�հ2:�6�⟸�%��J�-�*u��`%�lb>����ڕ��6�	sԛ�����mC�	�!�3a����:�)��UY�ŋ�3N��,�.2��$�|}������Bk�I�3�$���_�ݽ)�������9�`��Jd<�aB~Xki�Q��ܥ�t9�n ��6�N gCx.����}Qane�3�?��iVu�m[��tR ��d4]�ϲ���^!}��R�C�Ӟ�̎'R��#
�A�%E���h�h��� ���[X��$�ĥ��A��\e}�gh~�1.^�R���@
�P��e�V�4� �#HX� PiOJ.�&��'�q~> �SL࿟{��2�sԘ�VV+�IM�tҷ�1�/<���;\-���h�?�ؘt۩"��>�	ji�d����� �F]���hSH���r,0�^-�	ħşʰ���~�
6Oi���Ď+��5���۟����,h	>鉦�ԅp����#l�B>�2��U#�_ЛiĒ�+�̊J,�,��Z��D��D'Ī��*64���Ȟ�`>o�n��'s�zC�ƴ\S ��k���`ĬP`� W���@���653>�E���q�"mD�����/+��pĬ�M�¾Zk�_���Li��4u uF��z^�/�1�5�5�Nc���9����R��\�F��8���2T����2O���Ъ�0~�-\�׼��i|_�$I��?��;�0�(�U�}�*�L�W>���?*�p�����0:/Q�&��Þ����@k��o�#g��ag4~��D���A�RȨB�r^�V-��푵�A�"���"N�]#���A_�=�����rU7���AG��gw�at��C�Ɛɓ�������>+� �H�������Q�o��3��eiԞ��y'{�e�f{5W\h����c��,%F>�5�/���ś"\���-�S�Li嶅?ǔ'\}^�^�ay��\1�f~E��:�ku�>�o��!��dE�(��
� }���O���� -���$��O�~#�*J�18�|t�ڞ���J�[+��jK���e�v�I���N1�x��Q����y�2?�XQM��:�+����r/��E��-���_j��O�C���+���p�僂��я�������!�d�c����f��̺���X�+�0}멞�I���{�QBX^���6o�*��Z��A�@x.�,���t#DS!�+���A~j5�׻<�zHby���S��_Ƙ�"�l���=��5Ec�?TsY�	}did��j�m��9�xf�f{x}��(���n��{Ds�;�W�R%y�"[#:�.��k����d�4�4�р�����3A3�3ه��d��(���� ���a��"�����%'��ET�C!���9�`�T��[���d���|`���.%���5��/��pƞ�t�I�&b87H����Z�ֆƌ���ZksAЗU����K�.����j���o���)�T�U�$D��&j':��r��@�N�?�L=J��O�Sjo��Q�̛Yl��zVX4��+A��W9u������=���=Jy�?���U0��Q%�'�������� n��p�Jy(���T�7��E�dL5�,�R������W��81Ӌ���_8�t�/�zb6ϲ9PP��+$�<>y���?.���:9���0b�E�߸�O���ˇ��G)�߻V��6������E	WB����6`ͳ�>eP�A `Wh)l��p�X̮��X�sx-W�\9>2b^�~�Io;��������q����+���M���c��a�o*~y��TgH9�rX��ÎP���Lq�߫=�X�~�����x��"�ߩ�y]V�&���u�!�<�������R�R7&'r��˾Sk���d��G��A��x,��{��QBw%�i��i�&������Du�/K���V�
���0�"�a���Ŵ�gm�H�rN�=��/�D���	�W��%7���� ��8��zfU��O�>=��*"(�S�t;��
rA	���]O�����bY�Se��J�^�'.�ℽS&�R`�wu8+0v*��y�q���I@����HŤ�~��v�����S���Q׻?	�2yh!�;T(�?���-�Z�|G�]��SIەF����Q��j�&����ϫG�6ꐗC��L/P
�B��,���mf�bK���5�6����)�/Z��y*yT�N�b�O�� Rڥ�y���b;���p�a����e��k}6�)��0e�.h����s(�"�*Eg��5^1�?{�x�M�W�fJs�):��&-NjH#;�V\��ѻu�\jܹX0K0�]���)'�F.%f21��#�req˗F(_�r��8Zȶ���*�&�Aiۤʿ혞zSzS�]������:vHG���]���ls+47�mz��a�G�,��ڎ���w��6�9r�MB�yx&" ]f��,o`�i�8��x����j����pmO>��� 3%&|=���b��L*�$��=��b7�K�Yr�ZL����?����|���ʸ&�A�x7~���-��eqj�[!e��PI�4tK�D��c���-��m����u��[6��M�h��j�֢١o�hu�МL�KF�L`��9)p��̪�y/��Y�"�d���x�#�X)@e�<ȕ���o�y��B��*m'6&�/���<�U�(��w��D��eڐj�,+���X�D���f��^��iS�[�e�eҏ)��q<K;���4�lɢ؍<)�>1�_F��	�׈Կ��'���Ga��Zܬm�ua���<(���oaTX���0-��ͣ��*{��8N/1���Y1�xY��O���K�?��$�C�Ȥ��R V���z�/	���c��o��H��g��ˊ|�]
OL%I&�wy����PaH��S����G���J��IK�h��_01Af9����
�n��t5�:<�ģh�� 3``����`��^�q�Lѧd�`��DeO&�ZM�^�7>�G�k1β��9��'�_�Y�
$/'�@����]��BV�t`m��������Ĝ��O60�S�៉�+1�>�$"2��8��2Z\��Q]̍�/��);W�k�W�)��{��"ʸS鴈��ޒ$E �v»�Kmu���U��=B�۝��6���+QK�:�֠ �2�0���VD���[����N������,.�W�e��W��^��v1���S@�7`��ð0�qZ��Cp�����������n������ ��!B4b��K��P���ٌf��=�y�/�#�OqB	�|0z����!p�h�H<8��g*LV�oGӨ��ه���o�Ŋ�\��]zZ��Ȥ��@�ϧ��|�%Lb��y����V'*#t��5�����f�GS�ѕ�x��k����m���CdS�hm̀�6\3�B]Zs;�1���-�������|5��@.�ES�{I.@�pt-t�w�J\m&U%��Yd��1���c��lf��u{N��@�P�LG8�� $�J��H$��mZK;/72j�]S�e0��3A7���?��.T�����3Q}��	Sk�����E�-�����n��!��<�=I~�jN��|AIZN�����m��uY�xsA_��D$9
�~
�loo�K���jx�u��a�/��̑f�V����r!����s�EX��3�"�����
�=�/AzZ�a7���Ss�B ~���X
��R��m�j�2��Ϫ[Uuw�7�\�@���mP;ߦ���|3��)�a��]�xE� cI�tB�XJ0��A�pܧLN7���gŹ����Hbv+�����ݹ�)c��S5#D:Ը��wZ@��'�5V�}ڄ��ݵ|i�~�)84�f]%-I�)�q�V!�"}���[����Cǚ#���V�ͧ=�1K�TX�C%�"�n���E�j��ځ�/�E1׌�/<U��J!S�y�u���%Q'.*OFS9�����=����*�~>���c�qJ��P4|s}z*�(�L�9w�ֲr�<h��I���>�l:�t{�2��o��dj�����G�_>E�K���,B8��B��*�g�ͮu�Y��+�cdx�KS�a��ɵJ�)I�q�m���\��%��,��d2^0�M�������e�D`$E�a�i��u��0|{����\�ٞZQ���Mu�X0b�	�)��=A�޹3g��]I6���w��ٗя�_�
p�i3����s.:Y�w_p��W'C��v�*�"�;ݴ�\T��nq5�t9��<�)��bE������]~P���F4Z�\bߑ�����P�2v��%�- f	�+�qI.�m֛��`�wBN�bm>��0��N�&�Ņ�y��c]d��ь���Z�$|���p���Xc���5�+;H�c�Z�΃Ē*Tf�U�x�zԨ��L$��9h�")<�[����W��W� I����d����$OPz6t�֢����j�X�;plV�^�[��4D��^���~�z��$`*���[ȣ���
q}�G;�1��n�*�}��M�3}e~���B�(��'D�5M;zp��d�)�S<�G����D�J��	^Fs���*����0����(�/+|T힇���16j�ف�NP�)7B��⚓�`����st�� �C��!�ͫ����o����:�\B4'ٯ��Oo��Łj{)�£�+��[^�i���2jm�z�DQMXߪ���h����m��	e�ESMM���t�U$ǿ�|Tr������\i/^~�2�د�y��[��'�k�^�H�г$�̱�s��-_��^�Zػ�dL���RWR
�J���7m�\��eP��w|�T腁�u�ɮ���;2��	�7�祥c��U}c�&`@�j�!�x�ez �tg��H���a8$�ħ#ur?�1���C��͕a\���^��F3��10�پg�U�vʢ5��2�]��l��$���
#�����;�v$@!���u������ۃp�9x�&��&��	�:B�cr�Z��|o��)����i��hj%0t��i:`�Jp�|ŷ��~��H�ɺc0(�1��T�n��Nĵ�S��-j������v�c�$��l����N��*�Ȓvn$Lc�\������q��u�R3>�K�[V�e�އ�|��n�J������1�X�e���q�ߵ5%2��قZH]�^-��6D)�ң����ь��5��F����L�̮��c`W��*<���rR���a:Q�C���� Xvk^v�`rH.������Q��7�����^u�>��޷@��=�u�hT�
��,������F��)W;�ם���B�IMӖ�&�B*v��z;9���X��ϣT+�Cv��\�6���������>�ܖ��oΕ3��V�����o�TG���<s�Y�`�B�U]s�k��f]V(�򌆮w�<�٤��r��rX�dw+��<L�@N}���+E�p��N?:zK��� ZC����{?�!zxZM��`y�Q臈��3<y�x.�]K�Ǹ�"@<ި�U�];�Y&�J�t��
� �N�jM��+vݓ���S�m�܁09`��B&UV��G�D��M׉��Fz���)�Gy?GB� �Ŗ�x�1agE'����Tl�Z@%���<ot��z{�V�����O��3�qsN�蘜�(w��J	�S�7�H����}.�Wr����4q�1J�|r��o8�{;�x5��״Ϛ��GN(s����~�;�h��	h�E�!z�������?*]�����Wb��%�F#�Tz��
�
dMFү޵���q��^��0��]�.^�u0�!#�u;'���R����q�FzVcTɠ��R��s�E/d��?R=0���=���F�1��A���S���y��D(���&���$mP���`�Q2��3A���?���Z�02�Y9pF��tjݎ+�H�l�4�0�;����X;�_3�&I��v�;� %�I��So�]e�HĆQ�)����_=��41T�x��4�tD��8M�#Unrܯ&*�)y�*�!T���d����;�i�ϔt��-��)��C��*
֏P*�-j_xE:�x|<��� �,��l����pĻݫ����fE˵g/BD����Ȱi�S�4���]� �4Τ��,��w
v�5���w/���s��:�
��O�B	��0랷����S�a�IWG<&����6wè�r_�Ą�Q��g��4&�I'�FJ�`��Z�O����SIB��@��=Y�'KL��S��)gM��ݚ����;e7�2V9�-8HKwe��,^�����2��:��)L��ZX�[��2F3LArB#����[)�#����;k�	���#H[{�>�)�o�� /+ȇ*L��Xp��_B=>z�n�j��3h���癐Q�Ie��HU�`a)/*�3�_�5P���ka?����1E"��	�J�={��W�'}�W�P�ă,p��4����.��c��1u�G�6���rrE�"rr�[��F�;
�-��{0&#����x�	+n���6y���
�Jw?�[�G�1:���Ǭ�ux;.UTf��s��S�o��6�x���LF��2�Z�~�6��=´��7 ����\/Ѩ���o��ξ�[F1���ҥc<R�4�]H�E�jX�{�H��JkA[�%���Մ��k��Z��� 8&�A1�t�{���_��h��~#s�GF_�D.�w�M�J"�
Z\�6�u�O�x0Ak��c��Z�E<^f�~
ꨳ�ʼ��|壭��"Ӥ�u�]8	;����BGуĽ���t���}�&\�����7�[�g���Āa��;FNUⵟ�N�^�G��L����M�o� Wۏ蛫���&?�s�(��'w��\�e�24>�<�i	�#��j��B�����;H 'x0�D�}�_��9QLS	��1h��~"����Y��k�M{���EO�{Mu���/��"�(��i��d>H��O9P�DMѵ�wE�n�nB�x	���gt��?KNB@2��uc��ڢݸޮE)7��kd�l�mM�.������/���8� Z��a�K��e��iceǙ-�2�צ+��~g*�EdY>Q����վ���k9Uh�J �a��^�Ymn&�{���R��Rljʧ���A�g�0�6�x�@�#�o+�L���PR���PV7�i®������ �s��3ZVz�%!6��b)j-���1��t�ر7���8��s��Gr	w��k9&�f�EIz�]��Rg�,�t-�f@�u�GU�k�)7 j��iBºA�M6��?$'{y �p��Ri��!X�����Y�����s��o�*�|<�~	pg
��/�����5���A��Y���|��l ���_F��_U:����z����<��̽kO���G�%�t�s����,�<:zk���Br94,�\~;WB�.��pKH�[�}�Mp�6��]hǆB_�;x��[ .P��_���ъ�q©�K�斏E`w��	�u1먛x�UU]��sLYEKڠ��XKj�bF�)k��w�YČ�o�d}m�5�&5�'���x��=I
R6����S�>6}�vjr T�78Umy`��ph��%�f�9ي}��x1õK�#Ӊ�T�C<��I(9���o�t�h����'�YEd�EJ0���zS��iݾ�D����Ls���ق���%��۔�^�({b���SDa4z��0s���Ǫ/#5.R������hmOYVY*|�/�Y�]��������C�`e�ʾ��%<�m�.ZU��ۊ��B��n�T��0��W��+oD�8�o!��E:��|�P��$0B�o
6���|�-wu��.�,_����L92P��b�$L*O�y-�dǵ�ϚI�yP���Bc�O�L�	�(��Ϣ���!3/��
�ģv�m�@��.���!ԱĒ5E�1y.Ousӄ"�)��������gD�D�/��(�<q��H?��::U��#�Q��H�a�
&H���1���*��O��Z��"j_��p&����?�ّ�0��1��v�{�N��w[����ӯ\4��ڮS3GZUf%�l���	��Bcfn�k����	�L���G#����eZ�@��Q
@E(u>,�M�0�6�a�X�ݷ�fa!�r��|����+w��Wx��I��v�F+3��.�.��]�p���+�<�ƫ�Zɜ7���1?�>Di�V�؜A��pY�,������0-.��ִ`�'-��4�%�|��q@w�>.�S�����N�������A�3�^w�2����Af93/�]�cԿʯ\�8��� 1����u������bo�,�oR�綛|]U���3��Q�q��Q
��2 �&���3
!��k��p�����]]H�cI=�h��hJ��#*"�ȅiyͳ�1�\��Pl�<DF�!��Rd���@_%�]�R�&����#8^1���F t���G;Qw��K�&�Р@#��,���_�ru�)�C���H1��ـ�t�gB�{�м�+��.��:M�X�L���'��������R�hrs���\.I-��wn6������_
\e���UI�&T�0 ����'#��j��NRkX�KIU�)I&~$��ϻ;a���&�x�$;Kc.�u�A՗�'��S����Hx�%�?Ur�HA��_�<qS	ŭ��A�A�qJ�y�l����5GU�
%,�J�Ge����@\��~R�����~�4���ZQ�3�8_
����1c�C��)F���@��b9�;��j$���˶,���_����4�v�Z�3�q�w�I�n.��ê+������6�B}J����&y�ۊq-_��첈�N�銄��s��9w@dQ\�X[P���4߶6`吾�S;G��Q���$��ܲ�&/��/(�-�)V:a�A)���>�4B@Uk���H.�g�P7�,���n�+�h!��Z;P�(��$P�%'h��+�����!M`;`qw��V��K�:�ΐ5k�r�Z�����&�.F(PBdu�J���gsod4lX��nc9� �nұ�%$D��L�o�.���ye;�.���+9B�g�7ӕ��Acx����%c�m"��;h�P�t�0p��z��W��T�;=T�C�:�4�5}`4E�hQS�M��-qG�FB��,}.,O�vH���%~Ɣ������=�'uXͲ��)�Hq��~�:xd7��u�C��U�\��	!`����\�1����ZP�bݪf�9e�t��<r�>Y�1��B�-Nf`��|Gj?v┬݂f=�fQټE�����Ǧ�� @��1��O�P�޿4���yd�!�V:��u��U��(�#g��9��~~4^��������"J�w�ُ�~Q 1�dg~=*&I�RV�@�P�c����~�]/��R�,E����EϪ�Jm{�*G���n����y��/s���V�U`K�e�ń(,F��"
����dS�Ϫ��ѸY�n�e��S����HHBr�j�o(��L��q��x�{j�q3yg4��p.:eq*��;{m���hK��A�Ĕ ;ۚ���h#3��Yz_)Y�3SC������_P��������42�y�R�������t�\��]��h�(����5ӫ�u�Z�����
��+�� ��Voϲ5dX_d}���Ҥ��;[��k	�,�.b/2l�&��:�]|M#��X-8��$Jn����4ί�����}�����mF V�s��}�u�C����9������֫���2�^8&��g�*x_�@�1��$�� �v���-As�h��6H7"���eI���*E�
�D[Ƹ0�e�=��c�|+�hR���pA���3��u�B�{,k�WR���#զ�o,�w�l��x� >*J�el��X��������Ux���Ój�Iơ$�s���-��B>1��c�~�k2�E��T�Ȉg��X�r.�����%=����d┨�S�Hh��Ͽ�T�fY%�<�;�Q-�����ѴV�ۙش ��% ���M�Ku�Oܜ�\�,��������mDH�F#���w(7A���!�mM�rH���x�V�v��4aAUpu���	�������*=���Wߜ.��HNB�׆�r}y)ݜzȎ�N���BN;#"��Y&k�=,F]�7?eR�6e���:���d�bm�X�˰U�_����M�n�8�L�uB�+�ƀ����:��%=׾�͍O�߁"5���Ri�0j�lQ�?�{��Sjs�*Gr�����/����xҶ2/+�,������C.#���k�Tn�7���h�n4V��6;��oRV��ۑ�Z��ѻC��4�P�{�����c���?v)�{�_���]����R�ѯЊ��2���9�ܟ����|�H�P�F��j`�J��F��l
tX�錢X	��x�$'�t.�7�r`���k��:�r,�.:f��N�b�O��BZ��2�5&���*Ư�ؑ��?
0��g:���ԯJ�m�%/��4��;����e�����ԙs!�C`�f��
��{cV����Z���.�z�͉�Φ��S�Z�B�,ƉI U���+�Ehu��c(&������R<Y���N]0�4D�7��f;��o����0r�<L$7fz�����1�iΈ��j�b
�������m��q�����k��zF��Zh�U�?����ŀ%���f,c$O�d6�`Q�齃c:bp^L0d��ؗ
����.���(jD�f>P{
#���xƍ�P���>���X���������(DM(H"��c��@�,���-��	��c�t��+�e����<~�Ғ�}E��%Qx��$��dkf�v�S��`-��P#��o<+���GO9~D���K6řm�����,w��PNFmY�����j�&�N�:۩9��d����5�K*:%�J�S�b�	m���?�.�������˕�w[BPS��F���X� ��M�SACv�_^��S�������2���za����?��)�GCD��H<_�Y/5j$�������:��^���wp�*�C��!ZI���g�+�f\�/YQ=j�� L��y__���dݻ�HE�\��G]b=��� P|��e<�!��a�_����1\l0�ąZ��-^=t�,�L�ʷ��YAT�e�s�:��X�E3/���7�&ɭ�����CL&-��X�P�́m.���T�J��ȧ�w=�j�m�]H�#�\����2�ێ����������C�=*vOU5}�h/����;���8�X�ciݘ<�ƾG~���}���'��`�[k�}}��<��{���=k�:�6\���'���D[��5C�9N�
bQ������g���	'��g��QfL�,㦃ͨ�Ĕ�f�wp���ɗ]�4@�:6fMwR�����J����n�����T��q���O���N��qsD<qOk7�$���$������p��p��?�%��$m_eW�:n����Sׯ�H�]��-)M�Õ�&�e&������D�?QF���\�o�+���A�F3�Vx�}}U�x��w9Diu���q'�e�]^\Ŷ[	w�+�;��;G.�'iQ�|�[�߷[���y�i��z����)�����%R���K�7����z���ng��+A9)9�7���O)��|���z:����b�)��,��-hQIzח�p��OTSk�x)�^��Ɩ��S���8|�&�
Ff퉃N9��@͵6��>�}e���@'P��e*E	g+��M�<���g�*\��"�k�U�jWoIIU?s�n%K�ia����/Z��>t���g�%��!�6�S�~�U#؄\��?ƫ8^V�tq�Ol�Qi�(�Õ:p��ndk!/�(d��ݻq^�jT2����^��3��Q���5��Qy����͡���C��['����3���0�H��|�\Zo��;v����p��U�~?�5x��.�%{z���H[ ��@ �\ne� ̮!�[���5Uib))q�ցTk�L�V� �u��}J;�a�'J���ぬ�Y׆S�ӆ�D�O��:��s�;��O�4j�$5�g1ɀ�P�(�K]�~�7 ����4�-�L{p��)Ee ��j�"�6�����i����Z��ɀ+�n���˅��6ұ��Â_���j�m�U��(î�bo�̪�}ՏΡ�d�{�{H)�����O9H�c��D�?�j���om�K�),�^7g�`Ɍ���Ý��e�t1-!F�2�].�W�}3�6L�P���V�cc4m�b,���ܫ]�3��S�z�h�nF�����9���Z�:��AB}�:.@��Y�
Z�_�8Vb�?�Lqx�u8�_�����=`�~�ʏ�5iv(�hZ����h�S�p��BUG�J�*�6�yy��
�/FS�>�}߀�1Pu���:��Ap������!-���w�q]�8%���,���g
�.�����uT�#/-����C
��N����jN��&�J��[��X�t��WE��h�I���o"W	�?9^pf����d���X?v��*�[2�ja9�5\�#�DG�k��~�������x�AZ��l�Q'C��]�'�\���8���K|I�ċ�49���y9Ed�X� s[����	���7����et��W��m\Bm�U#F�l,/�3��5������@�7λ*�����������m[�R�K����pY�ٌ7���y	>~@c4�F��
Lժ.Y��.4�*r��/�Mt<S���R�{����V/�N�y�U��Mkʹ�u'��qk]L{G���YP�)Q�Z����^��SPO����K7�x~S��>)K�	��d	^ʭ�GJ"�]��\�j5ڒ0}����As9����l9�V0��3³B���ǎ�60B�t]7��Y���B��=0�f[Q�K�xD�х�sE]4E�B��
�Q%)R!n�6=�E_�F�̦Ȩ��o�Gl�'���,S�t���d��{(f�7�Ƒ�r�|����R��黈�J�WC_�|U�PV���d�^9��@��-����@�r��/@8�zx_{� x��<�r.��m���a+BcD�t�m��p�j�1b`����dX!�؂S�/���ފ������L6�P�t���#Ҡ�Vh��d�ԥ#_pZ�"�[N��ya�Ew����~�}�ވvV�c_��hí��t]YD3�Lov-O��%R4�>b��;Q�?���Ζ�`�xd���m��
\�1��u�}:�j&�L�CB��C�9����"�_���n��ժ���U#'���T�����Cjb΃o�[����犸�v�$sx�5V:�\'剴yLR*����`��\��Q��k��������`��jg������dK��-��|J�X�+�~��QUM�Y1�{ʬJb E�Y������^u���{8	)K34���<Ƃ�Ke���ko1h �^��ȎЗ0I���o�z��R^��A^"�S�"&��6�����n)�q��R������O�����ܤJl���V9;����Y`/G��Qn77˯�\�w{|hb��=�g���Hݠ�Cg��[����٥�ЎRF�
�bA5��&�E��gE�����DK��:�1��:��ԌD +�!sp1'Cs;�Қ?[��k?9qn�Mv.$�i�i� ӵ���[�2t�S��X>�L���Xq��>��ᅇ�w�*�%l��^����!�z>`�ؼ5�[�N"�%��
��Q�(2m��4�a�e�em�1ucx����t@^9R`���Hj^�T����8j���#��4���]���_7k����f-Z�# �=�J9���9oW�:���1��[�6l����E��8�2>�3��A���ʜXgk�����|�V�m����|���Ϯ�e1gA�@�l4��Mū��&��~�Ez�e;�2�H$�]tk|�*"���Q�5m��/%�k�Z<v�S�O�
 ɚ|����e�Iky/�PD�W�����t���W�:���d����M\�f{��<ϱ��$�X&^Bd�n�+�{A���o�����0���U$�W���%�۾�2��r���v�����#���2�[9�>q])��+�"��O��m<z���:վ���`�wR�m|�a��Q.Us���Rʬ��fe���H���riL��A��;b�!hR�ܥ�<��Ad���̢�f�lh���в���!tc�%.+_�E�4Dˏ�[SWCY&~:��+�����%��P�@v3���0�1
����P�	�#`�N4�ph�Dξ�{���G���Ф�/$2'Q��g�����1����d$y�=�cT	�e����@fS��(�GΦ��ɐ��S&�{��~co�K���!���Q�0�`kx�0Wz�旎`�w��Cc�e���o����.B�M��q�C
��,����4�b��:�4 Q~Ѿ4����/|�rXcJ����_��P��s`O^x�7qZ'��Xlo�fU$B��@N�n)�H@���Y�PG$Y=���Ot 4�dS���_:�b[Dʾ׳�7���7#�T�e���K�,�"�r��sCK��,RĦ˓��Cm��.���+��Z�v�����ݐ!a��@�Ң/��^j� [SB@��#f+��o����fp"Bw��5w��|�[�%��~��C)������6#N^|tl�������`� �`���1��ɇs��:�V�U$�����Ӣ>�ѣ��3G���P���e�=��'���9�D}�⤘�^(E� ���۝��5SD ��(1�*�ͥ� jڼѴ���}N�*��N����Ƅ*��#��q�Gݸ98V�D�G�|Tճ���)�)<L��v��0��V�����nzfFຯ��BW2],�gcG�{4Z*����v ��˒})���a�{i�_�ߺ?��%���^�jK���
�=Qe|�⃎��Ag_0p~��9�zɵSd�K� *�F�Ͷ�"=\{=���$_�c�T3@��.?W!�$1A��j��[!�xE{����ky�<?O��A��QRv0_~v��m��G��m�R/*�G;:G�	��aI�:HڬXk$�.��0�� [����8�@�7Xl���`9�a�fF�ZP�W�=y�"Ԯ�Y�X��ٱ5��^��T�\m�a_�{��زJ�v��(�0��&�_��D!�褳�~�I%Re�H	�8��W��s��kï��7���\�7��D��u%Z�h��R
GQm���5♙�ߧ#�����H�Σ!dup�G���j����v�#o_�̥�	�,���rLJn!��c`��&���
�T�	��tCs�c�{lL��|%��R>U 2�#���M��.G�z�$!$�m�3���.�+E�������}VԐ=� Q`�v�T��>�f�P�:},��*�A�܁y�7�N���5�N�}����S������H�S.x�����o�1g0�������1���L���$�K�2�i�(M�Hh�#NO���c���o�3a'-1l�>�%}M��N�]/I 9�����:IhJ��=;�����:	�����Ãڈ۹��Ԏ�G�I�b�&b�B#�)x�Dȷ1��_$�$��6y��A�	�dKe�ؒ��iQ��C�8�)�3>�$�!�b�;�%��~��2�z��R���Uhθ#�3�qi�$�j�$/<Lp`��;5��~�c���9Pc���Ұ��k��>_�y����_�_?c�ʩV���o�B�[�P��w��
��I���<��.�Lg :�Mx\r4�7x��LM$�8F#���%*��]	^"�vsl�_�`��Zb�4A�޷ɵWݳ~�Ϛ��:Lh��х��E��g��o�%]���<#��ɐLt3p��=W�S�q�E��s[��,����R�T�I?��/�����ϓ�y�����[�6[ ����F��������؉V?�I�yn�6���)���"��{jm-��Mݫlz��[(5�T�v�S<��q���2R��",�p�v��zx)|��O�b�uCs��	��5���6�� �0����%zg�����ے^����39�'�$)�w��y����vL3���8zp*�����1Wz���tU�x��x�Tq߼<�{,^���.�~�9hU[&3Q
WUs��� &^�H*�A-R1  ��;�'��b��{sP@��AϨ�؈BG��!y���A?2u_��l��-bʥ�V��F�kZgP޴����j�G.ĕ�R-�����Y�B�D�d�S	�<��$͎�OD̈!-$NN��YԘ��;�Vm��Ӧ�GEױ�P�����{�#��8^�������7,�붢�C�p���/�9���4i�v�af����t�jP�㼒i(砇������|��<�yW؆W�ʃ��)	YWoU���٩����2r�H�a�Zw#�M �Yi{���7��Oj9 W�L�{O�媿��X(h�s�oMB�Ai��o!j��:Ģ�dl$9�x/hc�{���)�rdD��i)-��������¸E�J��ZQ~Fأ��\� ��%YrGM�	��j��L�/+w Kkv�[�
�92hƣm$�U����*
��^�!Q�}�������00\�w}�-�1������N����u������~�iq�ゅSOP�奄�b#�(�q��0����/���q4R"���s#�Ƃf�v��!	I'<�;^��w ��ే4I�5��O��z�����ӊo�N�X�,��Dw�71�����a���(����Y��0�WE;�F3!��rN�m��j|�5gW��lx�$+�'����2�]�pzI0m��)���!�Ψ�~q�nq�*Q������C7%[5�i���ۜH�V�e�e0ɺ�N��$��9jݾ�n�`�mQ�� ���֧�:�,m#��%[�%���o����ap�/<D�!���ǓN��������Z΀E2�j9^ ��;��8�#٤.�6�Xk+��G�c2;@ɏ�e�s�)A���kFP���g߫�r/��L�����n�,(�BCF��I��ڦ%��{�P3F8�\�Hs�� �Oѕތ��uC�@{�uNgz�Ș���V@�.�IVb�������}7��I�q�Z��|Fg�de��ç�?�CqUV�c�0��$���\3I�<��m����Q� ��x\��xj��K�l��F �Y��{�<�������\p_�:�Pd�A��d��E��u��������:���F���j��^�����:x�j��R$�j)r���=)z���6���n���j7�b Г��";\���'�y˱)B��/��/�0H�0Vw�g0�~.��(�Q,hw�+�0�*s�!����JM�O�p�q۹�#��1`�B-'�x��PE��)F^J\��3&�K-�\��K׊L�>��6د2�۶�n�/I3���%,uۖ�yv�"v!�}3M\|�s�*�2;�m�z������Ź�	��r�P��r��O.�Wmc!z{�c����p=P	D��J�v�g]�XM��%�=�x>���g�w����`�=	�~F�5���;fa��ԉ�����U`J��I�����s�k�����-4�e��eT�I|cu���̿[��z�����0!r�5�-KX���.�����f�)���Т�}�R����Z���r!�"�b������~�cy:���>��,9��H�\���<�cd�9���]/���koo�s@14�5�ys����0���T���G�e�s×N�\������Y34��D�Cڊ�7�pg�s"F�P[	�J��<t�=���d��7-V#301k�����&�m�'jK��R/�f�F?��r������o�3ᒁ=����`\��8￧���6Aph넯2�p��WvP��ʠ�w��3dq�8���~�]pS�m�T�����m�+P��am�3ůLc{�#��bn����O->I^z6���e@�;N�1��a	�|c^j/8#�t:W�0S�����t�{?�Tw^���]Q�Rˢy�=���/l�����e7������r�'i`��u�R��|���:�sadL�B�T�e��Ɔ��NȻ4<),y�%��23j�Zq�s�����>AM�@軐*M�f��H�����*��O_��R�1('9ǯ��jN��6q��ϗ���uH@��Fk�r&�o`��Nh�iL��ȭj��/��z�����>�g̰rUŝ�j9��f�w9-��K��2��.�����u�1�E-Դ��C�Ѷ� ��Q��Rx�e�k�j =�v�v�1]n��@IŦa},�b���eϷ��g�#�/F�w��!Z�&��]}��xƝ�.Ӧ��P)�5Pz�2���a�����Ǒ�E0��Z����_X�����ݵB@�<��=���oM�3��pN��V�tF�&�TʁIA���[�8v���0�`-�$ԩ~�R��ю�a絬Q}�J��ߍI>�2���-���=�,�ѻ���Ztۃm�-D��d�cߞ{�I���o���6&�����+��?u��%�chez�J�6m�����-K���]��"�����l7\�p�tUԠ��>��IE��.梩��D��� }��SM '/�b,���A��? #=]�G�氹��ޚf��i��k<��Ģ��%Z'����d�[gZ*֚b�Y��Qp}��^�]�DΑ�W�C�ى-~��h	v�2�	u)'M�i��T;l��3�QO���B���o�SC������!7 �|c\��|������xv�֜�q1[�F{&{T��O�ۓH_��\08�����v6�W��mՃ{4����X^ĸ53�����}d�m�K�VOi|�\=I��Y��q��jnЖ���R�����Oi;>��W8#�V1��N(��e�
�އ�O�l�'��2��t*��b�d�+��2Q�ew�d�U���pM� �N�M���p�2��Q��?B"�1M�l��v���k� Ѱa���k7�lS�։cYϏ>tq�[���-i�Xy��ĺg �{��R��Ւʕ,2�LUrV{���_̖7|�Ը�F~K�Ngz�(�Zwފ3lW�ܧ	&�v&�n	6���d�9���!˵X��{]Q� �io����U����)��9u��:!���HI�n�AͷЅ�m(#�e�r��㇩�x�/
��f�R�A���)����o�����}e�ܒ��d��&����6��Z��z����z��s��9����u\���*�R�?����>��	<���*�/��,(B�mе���3����-]/A�~��9IV�d�$�gh���1������������VR4e"���k:3�~��t�7u>��*�WS�6��7z/�އ4�p����p@&)�x9Et+#��@�bQ�O%h�\+��#�鳏L�S��'�p����Is�Z�h��y��z����s7r���%ͱ[���aq�R%���,��q��ĚV���u�/ܜ�e�am|��9�/~T��rO�ɫ���B턯iB������۵9�Pa�_��A��a�w�鯓d�����r���}�[��j�U�ѻ���=��b��aO�S�N5ɡ"*���@�ϝ��6IIU"m�}������aN�>@���.�F��"R�^����:U��@+<��Ą�%���/oT�ʃƖ��cDH�A��gPI�����`9��cf��;ЫB��ҕ<>0q�>���o�� ʵ
��_��[g���
%���I��k�����y!h-3��HmA�G	��ő/���T&ep�	��T���Ri���Ӣ��[q;
�3�9v�8�me�7�܌�CEbZ�r��x�X�<W퍹��E�g���US_\q�ٍ�r\e[W"n�?�m��E*L�}/l��x����+�x1D��-ҕ��bJ�Cﶆh���E`�5YC��(���P�L��������-���@������
���泍m����^4�Wc��äЁ0*Z_�pho��L�[m��[��~в�z���q%�Ֆ�P�w���H��v��TOG% �+�I��t��F��b��B$�|�Pԡ��!��[�p{ܱ��L�
�����$Z��4g
��ѱ�g �X����Ѓ/�2G.`Zx�����<N��⮫R�G^�kxR�kx���B�H��ބ�vi*}EM�Ǐ�{����N�!H\9K��C��Ԇm{�2��dv=)/#�%��^@�'	���/I��\��҅�!m�?�&�%�]�!�a�[D�A��yr���X������N!OU�o�G��2�3�0�V�/�Da���%x47� -�R6uMO|��I�s�s�ޠ���`*L*�D�>+�_p �k�� M.8X�n�W�V{�9���X� \�ju���2ɮ��Z䶃n�XI�̸6����D8~7�)¢2��@DG�\r���w�Ab	��'�f���K����>�8��d���<�\�˧���<㏜3Fp�����T������Nl'�~��>9x@Zg]bB�QQ�Dٕ�(�ǪL��.�O�����^P~�	ɺ鐤���&tCx�}�&M�K�>S%6[�5S���u��y���)�tg�����/g����������I�b���� vr��Y$��:�.8������{�:�M!��\���UTu]qh����dc�18��e¶Y~t~*��pv.�
S�Jyʳ�|�qƩ��3Lʹ�+&m���?: ����7un�J(�B���bԕ�C֮Ѐ���C[��/Au�^�����_�҆i�ug�� �H��K%y���٠�$�ׅ� o�G|�dE��p5��c�����^�\��#6� )���Z��]��\���jVy~l �k���¤%���CzB�N�W����ZN��D(�g�F�'w��1Џdx���L����j<0����܎�y4�L�}�dFx�"?:$��e�W ��9�Y�s�ߘ����¶b�!)���.����
�B�D����Y�5>(@q0XE�{,���"���ڼ��2�E�UX��n�R@�ZT;}�V%�^�;�P�[9�0��>\�����"$������X��/�1P�����n�̻��,?�}�	�&>
ា��%�t ��j�����Q[��Ҭ~�<�w�%fo9�]B�[Y�W{�d�a7U�_������"�
� :��K��m:֦���[��KZ��6��J�k��7KB��D�<\��kь�ŪC� ��0!ӓ���g\�s� �I���9r��#⛹��՝ IM[�lVx��'!}!�����O�zS|�Z'��2��ɒ�C a7m�.[�;�>V��	2�x��XF��j�"�uӼI
W)x�!!.�\���j�r�߽x0�
}A^�m�
��{S��~q�����h�l���:����E���I�r��l"���0hb��'��{�`�߳<��,|
ْ`yrئ���M7g���N�jR˕)���ΫG��Nc�aqf[A�g�g"8P>��u�ð���[�U�i��� :��=tG�rq�r���$(�'���~Q,�)�����&��s�Ӏ��&F�(�`%y4�p�N��! f��u���}o@R��mM�ed*k\�L"�s��[��%[�X{|��)A!�fe���a��괳[3��*f�2i(t&�z j�<Y��O�����;�����Jl��C�Z���:}�I*oR�z�H2S��S^o�`���Py��4N-�}1���|�'f�{��^���i��
�)�}z
|�ц�=�z��n1�۩���� �˞�����L�n��L�ݏ�VF��d��dO� �KSU��k��g�+�d��"�#{��<v^ ��>�!�g�B������Xx�#�C�����Ig,��c�H�1rl��I��'
,��nI5򘥰Mdm����E{6��N�y�O��S{}�B�Ԣ�~L��9��\n��}���&�8Uw�5��Af��k,��!��N��Fru(l��a-�T2�#(Ȃ�]qK�E�o����>�ґо������]�]��'�F	8�%r��=����֗̬v灕>���5���!�=�i�~�AYo��5�ͺ��h�	4 ���ɽ�9w?9pmN����v!=�~U�=��NțJ��lxZ�w�I��ʹ׹��!�'I��u��Q�|��3�����"��e^I��O y]�7�=H/�r�J3٪8�Q ��\!b��7����	�;K,M3�(�'PJ�mW�w �")�_7H�ŏx�w{�}����� ��ڢ�c��?%�WK��=e�ř6P��0TA�Ԡ�Rlj��YEȳ�W�o`��P؅�Vˏ������a�������w&�b�2�/~3}�Q�S�Ʃ��Amxw�}Yj\�	~�>��L���O[=���/ϵ.!jΈk����u*HY�M�W^D�fq�M_��
���(༝Ѽ%�B�E�_&�γ~��M]�V�C��!��;�8�F�J/�[��W�A�6�{r��Zb|�á_aO�����*ؚ&7�Sw{�$qh�+�D�ʘ��mɣD�{N;}�+$�	�����(�]?m��B�.K����ؕ2�䍯�wm"���8����������5�v�JX���a����+鿬�����	�����v����Gwo5B{%�t�`l�����K6�C%�V,�3�R��Y�-���(��~b�����$��j.]�kI��н�\�2���fҿ�r�2J(�k죙�8���<� �P�ٽjcٗ��L`㯱�N�a���������H+�G��HsF�@�]��H�B!q�%� J,�PފT��l��h7JW�e���3�z�i�]����?^"}`�	�Hl�E3���(������M27W� (�RJintZ�Wvo�G6Tr��X)�����rlȻ	-���hm�� d s�3ӏ�D��rD
��3��N?�UZ���PI��& grM�}��W�_���Sh�a�.��&���3��læ��-k��T=��U��J��m��[I���� �G:uaR�!EX��5�;�n	�J�r�$~�U8ʗ�x���G �$T/iу:^�M��-D�tQAƄ%zNI-�K�h=E�D�v�Eۖ�-b�^$�?���!����]'8b��\39�K��[��;X���Fe�W�5�eP�I1V�B�_g����(���R]��i�G0�J������.�)/�'�����:��I�ԯ��y0�Q�:���Λ3^�����i��s�,�I���qi�tj�.'�T4`��P0|5v��o�d��`o����T���I�^�E�|��l�;��#&Du~ Yw�}��Ɂ���Xݵ݄"��ح|�o����l9O�cw�(�(h�U�x������shڭm��<�H|N��(�w�Ry�ٽJ	��H�@%�x�v>���QU��������࿄�̯q��ѡ�x��~�1��`�gF�=��ӋlO/ȓ�i,���'��c�b�m���$�m<z�y���\�I�_Rt��j-� R��X���JM�EM��-��N���֪>�)�*���ƒ~gJ���O��:
��\�{�$���q�L(B�@ #y��&�E�����I!h�ʡ����ډ��G���}���ld��h�w�?��> V��� ��t	�N¶�h{`D��{>Q4ϗ�8O�t���;Z��ys�|����MF��y_�U�����-f�VT<���q<F�h�k�1�Տ��]�1�"���)hC:�U��X;J˸�y��?�7X���4���P
� �ْ�C���jry2ZS,�$���!0@h�w���#�9���_�R@y��|��ib��`�������W+��Q��'�2�9iҍj���ڄB����28��L�,t�}�Bf��,��R�XeBs�WhJH[��E� ���P�Py���Iw����h⾩�[uZKK���4���y\�&.���p��e��hbs���؄�e��%��w��ӛa3KD��;���7���	�y�u�7۶�½�4�*�K���Ln�,��.yc��N�w����Ms�\�U�*���^.	�6[DBq_���Bj���2���t���F�M�eë<�j��uj�7&D��KI��2�1|P, ���Fg���#l�cdA����J��L�9��KFU<�˽3�I5?�|�F�-[���2S��|�U:nH>��'v�'�����I����*�_�ڃ�?W�9��8�P#t��G�ۦ�PtO
S��{��@��pg����N��ɼ���H��K.�dh�
#p�,��w�H�B���t��*kOk����8��9�a��/��֫C�^�TF� C��G�	br&f��p0uI�scM��!�Y�D�r>�R���1����`a|J\5�QN�z���7ԥ�c����<�"��S�ɧ�z[���	�S�[	�һ��N�t�W�uT� ���k |��~�s �NBD��/؊8p!�Ma�,��9d^�fJ���0j�{�>���-��� ��|�aD��%`B��T�6����k��a}�k�ރ���,�$��zu�� %m*U�[��A,~t������:`��MNF`qN��Ͼ��*ik�f����"W�������դve�U�����������m��@@磐>��9{�l&��]�L� q��N���B�awǷ>-�,�=�֤��>ދ�ݬ�Vh\�[ZJ��E8О��w]��WU��r�Z����@nN^��R咍�d��e^�iㆬ��n��"�7e��1������z)����>[d�|�
uyI��cv�t�>��%�G+�$d�
΋VH��X��{��;t�f�"o�@�q�3-�>�)� ��C�l��7j����U�]))�D��z�U��	���TЕ~�ٲ-��	�F&L\c��}����j5_[�K�E���C}4��ᷣ�[M����W�R�7�z�~�/6af����fx�`�x���ޓ&��QG&s쌍��e�/RD����F�QÀ����qћt�5֖���¬:�ħ���o�2U��Ӫ��ݗ7�4"�[�x�3DԋąH/G�SB�j`P�t���M��}�1�p�/�HR�D�5�y��N[����\�<RL�O�].;m޷�m����Pn��������w�]����|:){�A�U��*�l��[��3�;�<U�(�e�Zd?��o�p|���h.�H��憒�F��3����%�?ťԛV 7H�QfQ;n8�e��B��?���y[*-�q�]�7�tgfڅ���bp�'�Dٲ1.���+L��~,�.,��l�U8�����Sk0��Km���3B���}�*�d���4k'_�Ov��V;.�>0�����V
RJ�~M;�����% �o�֞=O��
#�d��+���#�г܉�Lt���F�1*�/�qt�y�X��G�G���oKTGe>i�*��	.��#&kfc���ΣSN6㯍�11Tv��r��Ӱ��3���Fx��y�� ��n؝d�ctm��>�ȃV]�6�q�LK���o�C����lx$@�0�j�N���R�3ݻ
�Xqt� ����3�|jrު��"�Q���d�v��J���_z���hx�F_��u��pc߮��Ȧ4_�0W�Xo�l'��n�5��H+1:�,y��	����p2h��y E��Ǟ��, y0u��V�Q���aR\	��n�+	��=�!.�Orb��KP�>��4Fwz�}=$�Fү�EU���I�i��|Whǫ@ W+1$��Kn+�ZJ�u�j��B��ʢR=��eS̽��Q%� OM���u�O�D�o}T���o1����8r����<}e��B��jQ�02�����ȹUO8��ql�-�ю�!{�_ms�0d��ؕ��.; �t����w��"d�����"�%ګ1�����1o֌؃�V�<��+�/0�~�����6�05*0F�uf����}������;<*4!Ց����E�BԚ�-���ŠO��2q;�U�iSN������@r��͔�$�:�"��̈y"�R^�v.H����� 4�*	�.mA*(�;�����˺y�_IH,+�P]<T�mU"�z�-1v���1<X֦��(�0-�_��aF����<\���c�*/O���,T���S�jj�Ҕ�C�U�T)P�Y��hO��&����l @�QxT�d�bC�^��S+֦�)U��/I��o�Hd��ݘ����b�ܗ�3!����Iý�@rr>���V9�8�s]�R,���o���k[hY�Ǟ^�k,|'�@�1�l ����u�|�v�2��9�P|��^���  ���m������X�1�X<PQ}j�Y:}6
<
Q�������\a~�IH	'Cbz��Z<�n}<�<�:��K�$�|��~i}ʂ����'�(4*�m �%��Ώ�u�B����/�+C��iOx����������̀,LU�I��}e�6?�{�^mv8NR]	ЪƇk��3��෴p�*m��S�ֈ�¿e����'4�Zv���������AaF��e���wV<��*���W��pW�l4����������`�$S�����"�����0=%�e�x���-8�Z��"m�_��nǓ3�i�џ�)ϗ�r-�+��'�ؕn�c(\o$+�xX;�e��dN��I�K��ucyY@�����n���~Y�DUX�B���WՂ�ւ#�}:^� �G�˖rT^�U�F-�z/�\���"��i}2�A�$��7ߙ��ʛ#	3���<��|X[�ia�7���b7�c�FeR��w��(��r�a��@��v�a�+OP0r�h�5[Y ��*؁�EW~�B�é�}�&N����R��wŐP��o�-��p�7c����ݢ��ı����W�����]��7�q��b-!���fj�2�+�Y<�Y�ژЊ��#��S��z�iA������#}`��^���&�C��{kDWM�X*�\BЉ&O����j�� ���ln�D(�x-�;�w���P�-"�KV�V:�i�z�V�	�1guf��o���:y�sF�&�Z{�@ܙGlC��V�)]�#s�ƴ	y������w.$�Ǵ]��l�b�bM\��a����b;��v�5�B��o�Z[��5Kƅ�j�է��pa�]'O��,�mֻ�FX*y�w��QN���>
����z��ZĮ��	�w��ZΡ.y��ϭ����E��9l��!"e����DPfC���0�=��wۇ�_/D�5�is��A�9�~uC�QY$I=[i��{\,�}ߪ���GgB�*N��o�� ƶU�1e����~���ZI���� ��u���UFǮc��Az|oi-fiL�����1v��:��R���j*:2�F�׵�N'm�Fy4��K���Po�s��&���%Ĭ�A��g���d,m��]���^���������.m����ˠ����2�+F��*��Lsމ+M����S!�{��Mq)��?��v	ɏ�ؙ��К��n�������F�Bm!�ϲҥ�C���X2����7'��\�\.�A��3��Lz�@�M-M���ϊ�7�ܷu��"��F�""Ȅ�oY�U��ogC&�9�8MU�r2�D�cfǗ4�2xzUY]��6����Y��Alzޚ���4#��y���v!��=�Áu�� ����(�
��X:���A�iT��g��i�t	B�Q�쁵��m��^X�t��9��� �P����IxJ��>��r ��9eI?�&���$�犯_�8^-5<�+��@�E�S1e�_��y7@B�X�~1�f�e�$��JP��o��*��N�p��)(mD��JR��(ݪ�9(f��E_j�to8�e�Yf�^�5o��YnD{<
,���
z��pJ��Fx��sC��C*L�w׾��FyZi����j4=L���]�P>om�*���Ô-��s�U������'�����c�Na�_��a�7���*g
�\���&������V׾3������E�,�X��;4��XO� �W�2�	��Z�A���r'�!��o*���1��Q)Be_�}��+�}YɤZ~�3�r�ݹ��Y2c������>��m�`k�VS���|��4RU\؃��I�%�Q�E;oX1A~�
$5�$�'�MoSʘFDo�����Z%g>p ��ĺR��vf�0��:���*�.�AXu�އ_�H��GӚ=�:W ���2�(g5�<��n�N��޻N�s���Di�������<��X��UfA�V����#�Y:f)�	�Z��Z���E��т�u��g�\/k,�_b�����4�����g:8*��=Z�7��H@��^eSq!�Ԇ��0���(�eH@7u��%?�?4c��ІگH��U3/��j��)h�mL�wu�2��Y�L�C_��sP(
��ʙK�����u����Ŧ���zu7�6^XVc0����sg�g.�L��%}*i�Y����֞�iD'����i��ȧ��ŵ�dO��'4�>�50EVCsAȷ�$�I�����W����j�����m;�~X9[��e�~ɖ��'�~ӅA��N8�+5����r��l�A|l߆W�!���;����R^���=Y	��sg����!�	�J��tZ�4`�~�����ThUK���jÛY���-�����:���A���8�;�?`�y)�`��Z����k.��l�k�;��}l{��>��v'�2���)G��c3xϟ�B Ѹ qM�Y����J�k+ ��r��F�{ ��B:S�6B0�!��`�>���d�*9r����D%fwI�Qz�N��	���aI�L�j�\�N��˕f��!�nN���I�{�&B�q��`�b?��&���V�}������#�Zҕ�$�W��6Y�HX���W��)�{�����w����ߘ��e[����1�_�d���q���2��<�_�"&��ͦ&[�����D�eR�o!a��]s��}�#3�Y97бFE�G5��Ϧ�"���s%!*�bA`N����V��ٶ�e}�&bń�]o�&Oci��I�n�ߖE<ǭ2�#5��a4]��������Ho�6{���t|��Y�P@�ep���+Ԃ���y��S�]�M)���z�!��7kV�G!ޢ"�u!p����Ͽ�ś��lG]�(��xE�R���ʥk�>h~c���~�i�?]�ű�?Βz�kE"��?㭿��
�;g|�chH�Ň����M���>���I��ԉ�/c���.s[�
g��|�U�Y �b��+�@���B6�)��.)�zJ��Wm�J��I��u�]�U�O��!�۰ĊI��&t���]4R�)���R1ɳ�¡���
O �u���)�Ρ��c}�����뒁'�����|�@�Lq����Ƿ��l���Ո�H�qq�h�qX��V`�2������~>1����p�etr��r� fG'u����Y��g�;oR#b�#��̠2g'W�|�-����+�R�h�9��+��ޥ�!���'�F�����cC.�f.��4���6-���-�@D���F���&Oy%�K�-8�U7<�n�o��g�7�ඔ(k�9Q�����/�W�=d�N�b��`/���EX{YA�^v��mz�u�u2���Km/~i���`T�M[g��O"eu��Q�
_� j�X1(����-�T��_#a�H�

&�N��[:�׫;0�$�16�K���-�O%�8	�>+��:�ϐ�՚����+u��F0ӎ����vEt`'�񑏡P2����	�u�]&s~�f�H,��E$�p���9�V��`���B�-i�A�x�M��jD�Ss]��Ր!b��i������n�i߿���/�����:�O���3`t`�������e8;a��t�<6�k�g�c|s��%��]hjT�R�.��rewA�R�r�����!F ;�j��ːrH�xF��cY�Q��FTR~A��6�+�+�f4�B��g�T�8
����[z�M��.h��g�f�"̥R��X�t6Cb�k
�P?�]��F΋���
�����1��~����$�����n ��<v��	|�xv,����4�xWI�dl�ۿM�bm����*�4T<XhI��2] ��&�Ө���sbO���Lxof�E|�۵o;E����J'�_�9�x�D�`$U�N���7G0�I�
����#�Գ��~��.�C���]�����x�E��)��?4&W�QwL�WųW���`^�r);g�T��[�E��s`�40��%��oXY����+6��j����h������r�ѩ�a|�E%R��@!�S|���w{%���n�5�O<}����]7C���j��a���P�0�''7`X	ò�^����R��/�����m\`{���3ܢC�n�2�~�9���<�vޖ�j^��YO���!u���W)Ȕn,$��\�B��Yп/!$*���޲ٍ8���hoAe�M2�|�@���f�L��U �����'�9��k+:b?���:'P5��<S��L�qe�-kd�D�#��+gH!MRm�|��1���e�#��)$���_6�P�p鯡ׁ�=A�}�U?9��x� �Y��O\�:�̤����]y���~t�����?5|`���^�z7d�ڪꀋ?�e�D@��oZG�}S��4`Ģ>JEg8ς����ؖ�mT�g=���!���aw��/��B#X��8�.�������>��\��!
���I�k{[ �
E�\����堢�_!("���hP)UC���8U���A�4P^�'��<��%K1 �4��������Eqp��ōx�#�<B������{U�~	<f)���n��#7�qe�/I��Ϛv��_�D�ޯ@h�O�f�t�Շ�k%�VSh9�	��h5�G�����/���j,CE�9��k�oT{�s2��7��F���ׅZ��Jr���f�ޕx�K�^�6Ҟ���E��7`E���ƕ��+l��c�a���@������S�'P����t�V��x]39R㪯�ܖ����|L��c|*�Bgz���Mn� �z��+g�P4�
K�;�	'\�i ��ԝ܇�ʴ��с3dY"4{�YZ��&y(긙��:�ҧy5��S�L[ύo�wA�e�����ST� 0]�(�c��t�DBA���s��f)�*Γ<v�6s&������l���������ٓ!$WX�
N�r�:����I����T�t��jT����?�qd�A$J	�d�R���0����2^/f�f\�c�t��*A�,��lHyT��?)J������nzT}4�eय़�K`�F�l���c�r>�t8릁]� �FꝘBk���T/
� �=
�dF;�Ʈ��E��f�㡄}	%KCf�q%;A9Cv-�dh-����Q9��7�z&W*P	v��7RBE7G��-j2;_� 	��9� ��7,#��Z�8e'-G�����#D�Sr���c�l���C:Zw������Ӏ�`f�K"5����1�L�F0~ 9�~�܅���QH ����2��Q	��}tܖr�֔�Pb��f[L�`��Ȅ���RY�:x�	��ڟP���1�'=E�ŞE��j-�f�� �����+�EZ�ɩ���n�	u���W�cȇ�d\_B�y|���f�B���܌��wWp�� Cl��U��M�ǫi:Mpx+꤯��.i�g4���%3�Ru�X�z�KP���A��k�U �rS��S��z]J[��U�M$���%5���5������K�K�$��\������9ص�9�9b�`��W[h����D=�g�j����"��s�#��[�u�K9�)}Jt��xK���|�D����z�גH�\��*iaW �k�k��!y�3"sU6Ɔ�֪����haK��XK3Yä��S��6�SuZ�� IB��`P�X��N��w�琓QI8��6#ryejw=p�k�\<���׼g���^�N��veQ� ?�����ٸ5����Hf��?L~�!6^sC��)�K� ��	�#R�Ɔ󚶸h���L��|�V�S�<�.|�p�L��L�&d5���x�ᆶ��{jm�q�$S�z�ܟ�=��;�=F 09 �7���^C�����f5�������ۣ�v�ă}mq�b,����Z�Ύ��Y5�Q�9��_Ml_E�cr�C��	%�qf۹���
NU�g-%�h�Kg� ���6p m>F���Zv���0iԜe5.�GcIF~[k�L�C \\n F>e�\��B��N�'ܜ}�P�#%�a�	 ����5P_�ܼ�-�	��e����rPl�O��D̙E�ESo�C�%ѢQ�*^I��W���,���6s�[�l����Hl�:��_����G�P	!rt��js5������z0�����|{�פr�G��xko���񃮖����iU;MO)x��^-'��iK-�N!G��9D����WO����é��Ё*���N%$n�,�u��+�/<	ًח�u�� ˻�gsM~�Q_�_�ܕ����Td�~U������k={��Ժ���	�lH3'��w��ː�k,�p�ε�H��3�@����)����y��2Q�y����kij�?�U~&�h��`�<*Z�f*�9����q�s�
�-�Da���b^�^��yj���]�I�t�7��<�Dh_�@w#Wd�%H�0��NɃ��y��5�{r앣�7��?x�vX���W�pS�)`|ea�;5D����x;
��J��,�S5�^�M%>O�-�w����,�`R�6U
d�߰�}��L�|o�K��IRbuY�|~�Gx�n*�R�x*=,mg�C��-K�d�_a���8ET��A�1e������y��LJ�b7�*�'*�yZ�@�乤_�y��-�Q�s{��ţ��X*��tZ8T&69!���@%)�0����ؓ4�L�dw�Vc]��#��y�|�	2+��PC��
���z3wf��X�f����$��Ź���E�p��-�p4䳿%�����1��!lvc� �Qlɰ$JlIK��d���wW�ۏ�c������Ygժ�CO?�U��@��OC�`�` �}��́6(^����3�FZ�x���N�:��n�N9��I�g��Q; �}�l�����RB�Z��8$��]7N�0͌�J�	cY;��=퍶@�U�Y���4��q���ܕ��;sX�^�+�¦m�h�H��~�6Po�Y�;[�c�2�%���Zsذ�<�#[�Ӗ,�N������({d�\�eM{��GŁ7��l5G�����A��Ǳ�(��d��!KS�2 �,MB8����>[5_�ury�C��'e�G�������\ǎ��h���({Fɲ"v*1�u^�6���_�Uy�����ro���#�Ry�K�ʔ9�H*�Y�l�iw��֎�ߜ����BT����Sy&b�O�;�0"�5�X8�y�u�I�ލ�G1cYxH����Q��MvV�M1ELg��Aꏄ@���.�u�n޷�U\�X������I��U�p�������]I.i�Iy-X��EDM!�d��q3#�z-k�> ��o\^~�p�(��X�e��av�@�������f�q�"X�k�1�Z>&V���w/U��l�,�wV�?�f�Q�_!�
,�C �����S��Ћ�r�y��a��2t����V��1�i�?��yu�]ht3��[�^y����u�Gy\|U�D��[{�I��d� �t;����kCMU���Ȋ��A>��&5�tB٢'���
�B̓���[���ئE�	�mq��Ro��z=G�,yș)�ul2/bᨌaKY,�`rʍOH��	�0؜���%�W	�4�Z1��g��!�ý��pS�H�q'\9P�I�="i+�x<��Ƙ��&V;�l%Լ�x����8��Tl;x2}	����d����8!'����15�����|�f�
䚏�Ƹp��9��p;��$�w�Mb�ѱ�ɏS���'/�];�x�����CB��{�����;�b�@��S{����ZQ��s�ZEO�;�Us����b��W�z.A�V��zhez��h�ݙhI�N��$����z�ٲ�=�q�`��? �խ4A�y���{LQ��:Q�rM���Qp&^���(�� L�B��dB�	�3-^�t(��
H}�2d����jj�ك��<*�ee,0��{��m�s*42�X����f���<�C��ut����f�/��N�#.2h�U�X�[�|&^��q$�JL�����hH)��[�\����a)g�#�3�?���jp��!GWU�4%��<���R�#(���;"��_,�I�F������vi�_��+����~�guW������/������X��Mᡋ�[��ɒ�Y
9A�
�Do��P�<�tV��O	� N��s�҈~��;���s���6�)�@H���;���^ �gY�iǳa˯��	v�Y�A��P�d�i�)q��#C|�Cp��S��y�8#��_q$��r�3�lWF�J2ݓ�&lZ_�?��`����~��y��^Tw����2�C�nn߹�˅�ne;Y)�ǻ	 �e���!�^:K[�r�nQ���3�2�Oa�i(�!QcGU7#���n>�/���<��m;��Ug�B�e@/����uQ�$q5�`��{8�U�m����X�7�i+�p�tk�|�&p�<үIsui̡�L�UX�Z��>�~-��d�O}�P�`�̗#�!�-ĳC5g�$��h�&��k��I����TmW���+��T�G�J	�@ǀYP������-^ B>,Շ)@�(Y`45��dl��D��v��M�n��*���� `$]�֨;�Q����}]�ܫq�ڎ`{_j�ǜ�J������dH+A^m�M�5(!QH��?�Hr�3x��lHl��>��L�Ų^omF��˼p&HT� �f���L<��ؾY!�!����I߈Y�YԩOL��� ���=VFRav:�˹;:`���$@c��u��'4�F�"�]����&G	�8(r�GϨ1}�ɮ�j=�C07/	�&6pP�/4q�a�k �z�V%� �	��a�k�*��ō����;��:t��\��X��E�k�Z�dk�Eal��2b>�y-��ɚ-�v�������i��h��@��!s���1���4i�:T��$k��Kx'��Ś�ƀO,��j�����emQ��/؇l���*�߷!c�5������`n�8R�N�.�;���V��0��O��Lz\*k����<`%�X�+�5�g��L$�⏞,s&�c= �!���
o�|O�ru$��s�Ւ�;N���e�L����;9����F+1ʮS��_j==E�Ԫ���7�%��dM��	��?Z0f8O\̵���̀F/�?�a~f}sfa�1к����{ei�	x���V=��A�t���;���l���vsB+�R.	J�kd����o�C����EE�EEN���섹�˅�a'{�cg=J4�>�Gq�S�K$v����v.rt^#�=YI��QY���!2��j�߃3��f2�m8�(2�ٸ��d����R�B\��Z
	�����r�{�Ԯ���\D���׉�גT�ȩ�B�r���̖95Q� ����ܘ'�efG ���3^�u�o��t48X0D"	٪,{����};��}�¥h���/83G����x��zQ��r��;���&m��p�钮FT��T��=���EQKe7��> ����l�Ƈ���@^b���<�p܉���R��M��VOUl��'`�%�7�T��j��/)��5 "��:TG��v�A=��ٕ���@Y3�T�衄;
�d�C�T?�[�𮬚6�	��}\u�T�9�0��_F��`Y�4�S���Q>�93�?��𲉮/�P�	e�-K��\�QE�<BusI�A({s��#5I=^A�_Gd��/���^Rڸz=�vw��rgU,C�xoT��!�� o%��!�;���]�I�����Uh �8{���C�P�@k�~W�#�-�Y	8ޢ���+s���߀wr�٩^�y�O���y����[�V�����e��C��৵�or���DEk9?�~ ��&�6ե�΄=�a0YI�e�|�w�~!�@9�	��Xʷ����@���_��`�vA�y����"0��(�rm$��SF�b0'��D��N������mpM�40�"�!��u��m�*'q�/�K�|��F6<k�J`T9��4_�6U�w�m��8M�yu�]:�a�V��\f����d>�	�	���T����9�6��Z����r�c�M�j����Ѩ�Ɲ�����&�S�2s�7P�����h��DF�! ^Ns�`�t^��(`��Gn���9ޏ���L��J�[�W��pSV�;��ϐ�	���z�L%}��>r�̵<4������d��u���Ro�SH�J8���	t4j���X�4��s��tg=�QB�H\�4��](�s������#|��Yh�����H�p]\M��K�ޕ�������f��c1�R%[�"�#������a��p[K��6H����ed��3�/�j��qe�V�_3X�T�D�C�¾�+�9>T~���٘�sS���i�Ss��"Iy�e��tY�}bv�伳����Y��B���9:t�X���c.dq�O�!�_���9@�$9�s���S�8'�\�Lj U����?���f��:����hcѰ(Φľj�E���$|ۜ�@HR��h�T�w{�d�8�/w���$�5b�=���˰���S����p�&�3���W�
�01�G�s�n�ܔT�w.2���:u/I���lR��d�{�����@�G���[T�#��+�#�Y�-�z���a���V)Wɟ�aF�`�;����@��M2$��i��E����cܱJ�8F�R�����F9P�p��i���E�ݯOԑ��S�O���	�ܚ"rb�]���ɘ��Qf�]�Ʀ��������'Ty��S�۲t@��@�
ҁӠe;WU�_��H�l�$g�8��	l:�>\��x����ύ�����Q�w��s�ԅc8���Gn?s+S�j�����߰�֒B��lf�Y�v7<p[XG��G�g׊iF%2�yN�N2+�5��ɲ��a�j;O����P�_�1�Y��,�n�D+c�_��wq�/9Hd��E��)�={5�h;X��}��c0��ԭ��m8�A,������v��!��n������w[�8�b���v��.���S1)75�u��+�0R\2g} C�ǧ������ %Y�O;�$��Q�c��^e�����[���e�ge�ެ�L�Q"�D{e������/N�7?�A�����6U�P�+Ϻ��D��@�E��ԎP�,�c�Οghna�2+-"�i���͔`�~��X]Ias瓴�kD]��P�DA���pA����C�DDet;�`��d[I�b<[�o�W9�ֿ{�Fq�Kk��/��^��x���u�|�����������e����Hf�VF*M��^��n�e��~Z�6���������AP�EP$j0����x]�|���� �d�$��/P�M���S�vo+��R����hh��6I�Or�Z���?`�;$��ED��}�j0�A7��k���<�$]�-�K#�����������]�Έ`u�)=kZ���X|����&[��%��^�0bV�[a1e]C�T0�����^�χ����H��ո��f(T�𱄪�
��t*�6�L8�Z� :��k�؟a��ƊΈҧ>t?�)t��UU��&\!�	�{@E�hMͲ��]�w?���ҳ��LdJ�f,�Ь��ϛ���2!�����#�?�Ȧ
�ey�>H�uO�-14۔"p�U1�*:v�,�AF1�@�i����-���<#֞�yc g/�P�廤H���^o(@�3�97NQCM;�|0m���Lk�w�d(W/*x�܂�2-��e/���4C�<��Z*h�όd�a��=��^>��%AS�F���G�m�E����\
k���|CK��Qq��0�	�������q��kR�t��1^�R���~.b�^5o��p��y2�0�� ������$������B�^�y^��ݨ+�}������].A�K���N7_c˼�����V"�>l`/v���h=�Nn���C�KxB�FQs����HW��I���ӪܛQ
F ��wgd�αc�r��p�AX�I���9۞�K�%�Þ�zh3Nxtx�|�d��Gew1�ο�g�tǙ6��u�^���kr�b{�Zy��j�I@���%�5��[,t���?�,?*�j�{DiK�&xZa�:8U\�4.Z髝!ļ6���+O�.�x�X
5;*w����y�s��L���"�|w)"�B+s�M����+2(�b����o���z`�T��4۷���q�Ɏ8����1F�J��ϲ�����<A�֚Tc�YC~#��zܰ҆$�,
3�j��V��������K,5u�|�x��c�m�+��_Z��ӱO�q^j���X[����^_���~�Ƹp�������`f4��s���4Z	�U]��Q���4n\v���]���r��2Z=muk� �F'��*.ff�
%��DU�(��e��+�JL�>ðq�2+O��%�y����ik=q�PA�܅����b�	e�gCɑ��]��8<A��(vA��y�%���W��4�W���n��$��:�L{��Z� � grM������YL8����׽� �Qi�>�T�����t����n�2z�۷�)ņ��c�6)�]\�Z�����oE�l�΂W|���?�5��^��of�~Z-"�^R�3j���= n8�Cv���+�&"��u�d�t|4�Ф���s�/K�'�8	L��Q�$&����Vګ�Xe��1|]	��~zC�������F����v���w
�L͘����A�'�s���#���-8��8�*�7B�<���
ʛT'�0A�?�5�h����m8Q�ʄ�n���n��^���:�s��4xg�v�m?KP @�7t�n������[x�X����@�NOXn(���9U�5�ʡvAσr����Q��Wv��M{X�1�}�Ś2g��7JiYl��KJo���y^�(�`��J�z��>�!a�ww?������:2�n��7��0ـ�(�UK��?�y�$�9��,1m����2���J3W`�W{	_�ڴ=��F=Ĝ1>D���=����	!�H�읲d������X$��̥>�l����\��pS�Y�����_�Qk�zV^��HQ�7���Pb�;|�2��-,���G��S�T��G��l�Z �۩��҅˧��"��BkVHsR�꩏��y(���{�b衢`��(�f�1e��yd�~M�6�T6t��*]��C('j�l�������a����3�U�敚Nr��e���shWz�1;u��Z�Q�����Y@�����WHU\ W�S��e#2�P�ޙ]
t��C-�i4�;��~:�8?��[�z����<~�����S�?`R ���+uG�!i$G��Ft�����
��/��)xqp�a�m��- �����P	�# ͅ�7����T�aԒ��naua�<DD5芭b(t�s/�y,��6�W@���0<1�>�?^#�/SN\��L`�[��9�.	���ۘ����۲:�{<�����
��l��o����k� �2n0h~\��"M��^����+����;��R�n�&����_E�J��-4س`���7sl?�%�G�v,�O5����_�ե�`����Uo�)J��3��C�{�����v1����ԇ���f��ak���Ro#r/��h��#X��0\�}7AUS���J�UR�
@�a���>��U�k'��
&7�)��
��g������:_�9�c������L�7��IgT�0�Sw`�l�|_����$#<��Mm�1s��w]��6�|�95>���m��'���*����GH¸R�����7�JB�;�Im����K���"��h�I�]V��/V��jD�ݴ��K���y���S}����[���C���9[�MI��"����É����<�Z.�~�=ǐiMg�T!oL�~f���]�l�#��i6����k$U���]�y51�Q�s�w��0k"���#��)cZ+"�M��S��P�O�o*�Em���/GsBn��՞s����3-�k��>F��-&w-ŝ��V�G(��mߜ��$c��)A�g��2
Wd���!�[6/�t .6.�^׾<�AKc�x(�$�Ɋn^}������`��r���dyq���c��j�J�����Fp����R�KګL��5`w�B���Sߞ]hpB�,���Z��h��ZA�-XTC�\���i1�)i�X��%�����]��>�$�� 6�ʳ���bsU"˃H
�K�ҵ'm"�Uwƭ�6`�g�Z%��>G��s�r)�+��@�DJ�܌�]�q,W��D9��5��?�%�3@X:U�2�
)ƌ�7_e�L���3eJ4�K߰��;�:Кf��/�;0�.�.�0�H��Nm�gE��$B��{��ft���~�Z_�����|��3j��3��[UX���P$�e}���H�Wd�*F��_�`��]a��و_Re_�.'pm��rE�`7��V��b�!h�)E Ώ�g�K2�U&(�R���18�w�f�,��N�B��g@�Z�D|�9�~h��.+�_ѐX��E�I9o�-I���MЖ��)���U�v��"�D�ך�^�k�
,�	T�
���m0v�؉u�����$-�U7� 	͑�U�?�5����	�Uh>t�3�2���^`�cw���p�_�YEO?yg�Ň��s��!M�i$.#�?��אָ����kZ?9;H�JyŊ�?� ��Ȃ\�]�:~5�W�wK(�L3̷�Al��E�_����<�w�/ ��1�{Du��Ƣ+:���S/�6�X�F���M��cC�pQ�Åx���Fu0�Y)Ε9̜v�W0G?�=t�6���U�(Un+�g"��M�%���L�A��h��x�9o#�]���oo��t�)a���8�г�3=��b���
}�px�Ą<�w��t��4��ߋ�2��}�Mt��-z'r�i �M���1�pM�C)iڱj=�L���i���]�*~��V�2�0�Z�NNX`B�,x&�&�D���_������B�>~�~ZH*2%ck����I��k}���G9\P=2�6��.�}���G^���� 9��!'z��Z�ȾV��X2�L�9���0�v�dgW����U@F{��S$ٴx�JٌYX�e�ډ�<�Dҟ�QG�PR"zB���m �,1E��Ju�zif~Ē��q�=д
n8�>�qm��.m���
 �Z��뢾�#�	1�v9;��X�����A���QC�eɲ��w��t�Q\n�j0�C���j�M�a=w�������W���tݣ�k�`Zz����A�#_�P>��ϰV���Z�|ϗ�DB?m?��͑wP~x�������֚��Q��q2�f\�Hi��Y�r�T��p��&��b�8q����e��A�1h�o��+��)c]�M��(�H@e�[��#4��	 ����� 9拓<����V� ��9�ɪ��R��,�6MF�Qm�ɻ������Rc����$� K/O�I���p���l��� O�j�崠�׊�Q�^s�@��<fZj��Έ�e9��ױ�g��܄�>]�n��xZ��YrM8!�&IVr���_��������IoS����]������9��I���S�Ԟ�2��Lt����06@q�A��GZ�Ft/�Ac�W�q`��i���:��hE�xY��>�4�qD��#��%�]n��=>V���n+F.R;޼�L��h�|��.!�(ͭ�0����^ȓG��Kב7��������H����\
��Ο�!���QL\���m��������i�(`[xI���+v��n��x�#�J_�`���j�t��
˕�s_n�E�($�>�N�[���|i����x������:}�f/���3Bc8�?��Csj��#8�vmJ�bWQ�p�&�VE������X]��`յ�t	���*�k=���=	u�ʐ��9;���f-4�]Ǽ?lX���6.]z�,����J]HS�2՝�O�@�*�������RT��$Ԉf�;��W	�ڞz�c�O2.'4e�H��[�άQSGu�ȫ��V_E��ǲ����B�]�Y|�E�CYU��nb;ˊ����|��SNl��"9*W�:�ߙҘ���l���~��Ctҷ�HF�HON�`�ڨ¶aJ������	�ԓ�_~ۿ�r4��-;�"��z����gQ��gU���'=ڣ~�5|�2fҰҝ)GDLxWQ߯��Ú# ����������&>}s�`�]�� ��_vը�Ԝ���5W2���ڟ�A%�4�_,@|a�}Oh�	/�`Wgr�͌�f���
�q`Q\���
��awA�x�l��@�v<�ױ���T�Ys���Ej'�E
2�1�"F�8�T�at.�lѲ���VZA2U���'Y,^=-�4���Mz%b�ωך=�OV'��q1D�vf�h&[�`�Bf�����pN�K���]����)�n��L�e]{�^g@��,��I�U��1�M��w,'e�3��!a�qvm�X������Ɋ/l�r�uNyr���el��XBo��I�D�����e�Z�#+�:T|[��)Q6*�t4�+��: t˛~J:�z��y�2T�o��u�����P��KK��pl��?5�Ĥ.-�����i���a���啨c�.�6�b#ou��D QБ�I����+��솉,���[���'_8Wv�a��� g�s9D��F����0kW���b(�#��w]\"S�]�֡���n�d(�Ғc]u
�Y�$3q�����}���K��
v�2��Q_桁��g���H���;�(��#*	�03��&nn�c�l��/�[�/C^
���	2.C�%�Yn�����x������[�\FD��fk�_�@|��A��Ő�z'�{�A �i'7Z�#>ʳ�%䧵� )�6c���Nr�g1����]+L�r5�˫=�%�#���R@�������	�Y�(?�z^�}��z��~2�
�Y\9�l ��d�AP]��Q� >3��I�}?2_(H��t��۩'{�䚒J�����QӚ�u�ƠRӋyz	m<�1}�*Q$��3��� T7�lR��֎�M;Ȇ�#�	������K��\/���7 �#S [�mO���S��;�!+Ufύ��M��i�b�c?Qu)��qa��z����wNŐJ�������+��]�p���X��Yl�9����|P�����g,WRQe�ꇑ�R[�S��!�O����nʏ�<��p�r���Z?��$�f���*0�!R%%r�D����yK0��+�*�=�V���Kqw$Et�rOa�
�_�ڰ������6X�&K����cޝ� �B�B3\�q�m�8���]����S�fA{�p��A�,;
�s�i�[�cxG+tۍ�	���+�fd��H^
1�4��G�Ȫs���x�SL�z�3�����N��oBk�@]��]i�o�8�������x�g�طy��r��*.팽����U@��U�Pw�¿�ҏ�k˺�Fg�N�@N{{2�v����&U
؈*�[o8)�iBJ�!_�&�*sSǋ��΅"U�$wYq�x�i�a��H�u+���>�X�pO|+ޙ��&�Y��:�ܧDR�j����i��my/[�X�'��ܟ�v�bf}۷ ��W6s׫&��cV��uBJ�r�����)�.�����^Y?F/������Ǔ �
����H�����Z�-�(<,����%�j�N(���^��+ߠ��d�a��l�W�����Z��@�Z�d,�D��G�-B��@����!{=�m�%��6Q����j�/8�p�o�S�������Z�O	�+��2}�k �ܯv�<E����R!GK�h'x�}Cii6�O�*��V���R�q���
�i'_Of�un�1X����KxPi��k�N�Ac�%D��㬻c�5�%,��v���i����g�[�P�7E����2ٓ5o�Zv�N�Z��E�)���'
(154;�>��3��Я�t#[�4�b���R���xUr��]�F0�O�뜔��B:I7"\�
؂8b�EГQ��£�>q�����Q����!����F�W������]ȢҮa�%�N,D����&�� r��H���Й��:��0�*/l��۞�P���i^'�T������	op7�hx[lP�u�>v��O��rQ@#���/���Ǐ��U
8�N��)�K$q���<8̿��X��*�BWQ7i��o�&���!��p�������[��b�W~�Ɲm6k�d��VH:)�0�i�՚�-p�=퇍kU.����MnU�|�%��lOC��L2S�����L@����S�`��}	 �:�ד��:���ߡX�,ȧ~µCGǏ`gۿ;��(ܩ�'�Z�/S}��K mv���8��� S��	됾ň�m{'�{��f[�j��/����1z3<��]Ww�m	Fj��P��o��6���ٿ\G����)��^Sh}PV|�6*'�>�V��,#!��}�QzX�낽I��lPu��\A_/�h�D�_dBf���m������ڐ�s��`��$�7B�\�dS���F�z�.Q�EE��L���A�����XOa��xI��?f�Ѐ���Q
'�ކ�����lZG4�)40�i�^ŸCb���I�:���VbL�@v5M��ѫ�>4B>�E5m=�y��;
{��. U�\r��л���fv~�a/��.o���Q�t�!V��������q�������%ښ�LPr�;^�0'yrgd�KPo��ÒzPi��ɯ6haJ�bj<fTf�\ ���#�h�� :����\{�N@��Y���=?�n�@>Lӣ�aj0�wXƙlH@�v	�����������j&�8kV�·8V�gd�ߏt�?�M�A�ԥ����Ǩ��_��eXyŏ"�r 
���.�T��	`��G�~0��[��H��'�qH�a;�	�d� �o>�N;]�9&}z�e�*�r����s)�\�.+�̈́w������0
p�� ��B�X �PPs��Ai ��1��i��a�a�v�����;�Y���9yO���'gά8P�/a\w�d�Ҥh��q�E[lUJ��e69���=�'�5�6���>� �m������9?���lJ3���n�[
(pBq��4s��B�O�%5������U���lC��K5�y�e�	�*�?�N��⸡]v~/��H�;Er`1�ue	�V�K9���l���	�5Ǌ�	�(��i����F�����z��
=��G
mRL�1�<"bn͐s:��g1/�4�5tMlI>֊���@G�'ؿ�r#�g�4�I�V�h�c����,�-�, �2��G��xL_�B�Z<�M��d�T��WzU���}# ҁ��9ga�K��Hw+���.u3��ݷ4�dz���/�i����ܸSps��+[��f��j�M��ȑ�&�pC����u�c� ��n3�w쵼5���@!h偟afP>�UߗA��&Y�U:Ƃr{H!*É~p4��MI5\��`?�/�4���C�������?A�aO%�b��Soyd
�yb�F��M��Hn�P$d?��`����c�h�&��]CP�� AM�(V]*& ���5�W�ʥ__z����T��i>o�y���X��'�.���Km�-����6���_U�k���7LT�q� �~G�F��.�����q4�}�=��>I��u�Zx3�t�N�o�z�;ؼ)�T_D��w�X����9���ZzG�E8f��IkI0۞��,�{M��~3�7��.��
�46�
?��ku���kQ�����'�_OAek�	i������:
򪋬_��b�����tS��ArA���bu��BE1���1�,����^)8�ͭ��4)��U�ڦ�*��dfp�㷂��Lu�(�
/��{MUU͙�׾�~V���w�����j8V��eA�� ��TZ&N�G�:Ę���|~�-l@�mXYOH�
#E1_�;*{�(�5QR���}k�伔�� r/�`�X1������\�ɶ_�8��<B�C�Sy�a�S:��³#��7�q�
�N(�tƛk?�en���_o�r��|S��������T���ud��8(̒�A�D����d.��U� ��}aOy�|�V;�i4���P��L�F�=�I؇�^�dM�hP�,Ui��0�mdT8eFCIV�ǋ$��ety�1���^���mnQ�M�0\Uɸ�o����s���19�g��O��E��j�5���R�k%btQ)�Ϫ_�Wc#ČL��jNjTָF�BW!��M��`~%?���8����5Q��O�g�P���^1�KW|�V�1Y��ܸ�����r2���A�G:A*��ƽx|[�m.�fҨ�UEֆ�@#>'c�2)����Y_߬|�f������،�[޵<d�Q�$�Az�}�7m2>�~��� �EM��e��!4�n��[]T�I����n�bmUPb���w��n����ѻݧ�|�~� d�T����6�&���]\bJD~�jr-)��Nk�2�/��$&������c�oڮ�}��C��O98y�r�K�)v�"��t���D��B Y����6��� ��h�!��ǓK}�p;�y�UN`��r��.���D�~�7�L������f3�5ё9?��G�nۥ�5+�1|���۾�]V"�aF߮�[�s�6SK��Ć_�R�X�R,��"$�dqB/�*ue�@�������E�6<�+b�s���
�a;�
x���?�z��tЄP��zpJB�� ����S�W�3�P����z�2�x�ui�'�*�"��ճ�����t�ݏ�/�G�Y�J�Ig�q��T�Q��@�=�T��i o���
����`�p\�b �ڰ��U~b�ԯ��,p���	4�K&V3�ݥK^sQ�����cH����k���~O>M�.�a���;��)�q�+]�/ף>�O�� �P��F*�e=�ی�q՝*b	kYD}��R#�2qˏ�ބ��v�J��)��8��DoX�6ke��&*���/� b���0����V�|���`�a�;c��>�I9_$��%"��  �B��;�$�ɟu��gh�譔�ش��6m%8]\����?�q��Kƞ����xQ�r�k���q��z�B�ɽ�!�Y�3��k�@��r���i�����h��{y4[���@�f�&�ݹ��0L3`ỿ�Γpp�.�c���7p���dd��p�*�s�Q�@�Loiw]��Kd�!�|Fڪ��.4*E�!T��^���fE�!e�a�/���	~�TuxLq��~-hA�m�H�d��h���p�(J��Ԭ��
��fm�G�!4�ʋ_���:��6����ED��ق^�f3��NJ^��Q���uӥ���¥cC;]E��:8{�;=OÍ�<ެ2��n�͒�iX*IS���q� �2���8����M��	8�k����h��h�����6��/��Є���t�-+c����߫V{q��"����ݿBڰ�m��I�i�d�$Ƹ.�̅�.�����'=��2!���&(�@���|�Ɨ�ժ+j��ۓ�:&��#�++�fstWqX���&H_ܰ0�4q��3��8ES=���7P�O���������\���/�Y2��F�ɀ�A�?:��t�LQ�I�M�Ɛ'pB7JN�������]V�8i=a�2���ݻ�� 3�H��8��]�^��˛�P�~�����HF�Re<�iA-�|v�,7� =+N �r�>[�3�.��e��B�=#9��Y�h��nTܞ��WF9�~�4��z?Y�Ӣ��A(BF���rK�t"&��䐄��|�i�YY����$!�<R��wg�=�O���W�MtY�?�|�����!�풺U���I`�m�f�MZ�S"8mw8��n&&� ��^ܡG�s�������4p��p� �1����3�<��pU]���j U˶Q�ea�k��#W�\ȿ` ��aD!V��
s$L���\(#��):��y��������H ���.��Q�A��]fS��*�v�p��iE'�XlJp����/4z�P-'@�F8]�n�>*�� �ۙ:�x�Zt�/���R�27�#s��>i�o���H��Z�Vtt��8���g :��Ôrn�v�M���f���6���]H�rH?��H(��R���T���,k�Fq*�5.�U_+�G�,�Y�i��CT%�4�7��ވ��I7������i!֌�XT�!r��Ey��B��6�m_f�������8������T�k�iM]w��Չ�<�����TiI�c!�z���ٳRF��&O�,|Hr�]��us1lnB(�~vg�@�nO�l���W���{���bx,MK���s��U�
����'*kX�ׅ������z���1�_ҪN���%8R�פ���Q&��e�-^ �r�p�����B+ߥ��U�D$�Ȣ+��W7�%��|���͚0�)�����d��˾u(j�C��u�*��;�o��Rg�H���3�K��(A�3Fuq�\�2���\�`�w���b�q>��A#	��U����������B���GO��/`��T���h�g�a!d��C��u�*��DZX�6eڄ�L�i-�k����$Ѕ�IP�P"�7;4�1�<ʎ�(����z�y}*��,{��k22�Ќ����<�k@��,��5����:�jw�2�(>�Z��ya��X�$�SF J.�t�*�#f)�Ww$D6Л���[u	s>"NH�R;k*|_���cs����6FM��\������쓁u��_���K�կ�C9��?��w|{�k���t7�c^�"��Q��47�����aBq�8[�~H�ň��R8�k�.��\������6���X:�6������f�k~�w��&�<9ы�b���#H���?7�c��E�ԌVx��J��Z{ađ�J����k�ዿ ټ�b�'h( ��D;C{~����1������'e|�|��F;��<%��s!#����\c��a�����Бi��BU��iYPXar�B�?��WלA�d���c��v��-�y$0��R�5[���H�g�C�7E�X5���܏�!3�;S�7��:��?%hT{����q=�,!-��!��ɉ��K�:�-�x����7�a��.���!!p|�����қ,� ���{�~w��jw��s%��IJ�{Ն���x��C�#��X���o,j
�ǝ���h��O2�N�q�������F��cyXm^9�9,ĺc���
�0��Kt�`E�(<�LB�C̴\T�d����iP�5ѱ���RkQ���7���A|L�G�|rS"�JbR��%H�;��Fܡ�!a$�5��1h���A���mj�b�S
 �����:Md�����N��&�s;K�r!�3���!S�U�M�gIQ{�QZQb��t�?b�z�?�J�54�ަ9q|��^�^��
M�I>9��]\ �!W�c°7Xmj����ٲ�ɖ1��YKd'��X��~:o��<?�{�b�&6��[�ztY��rP�O��p��\WB#�n���g�Y '�`�����21`A�o�)}8��I�͝���B0��)�hI�NIӽW\�(��[�M0���;�}�"�w�D�M�iX�N����E���M��!���PX!�m%}� ���A2"y��[FjAF~�1�I�˿�jk�B#��}̙�F���c<������ӄ^���5�ќ��	����ȑ����R��pO;��AgCu�F�SQ�oЇ�*~b�6�k��9C4��1&=L=}z�r
+��"D��8�o���*ŮT<c����k�5���?��J��X1�;������Ψ���î��˼M��E���D��	�z����!�ځ7���Y��{�#�(v\��s�(��TzC��};����`�W�Z���x���1_(WIV�!������Pi���8O=^���u��ۓ�;3���SW@)��覽�����Tޘ?����GaaDzyVV�k�#�V�<'Q����N2��{��?���o����B�~�nk���D�Ů���ɾ��sC	�YzM�Һ|JK�*}�.i����gK��*��gžV�!;;	c��E���o�$�k}�SR+}� ^��� b2������gK���z>s��]��a�;zhBX�?1��\]��D)چe<7��[�� �
@.��m<�#F�֕��]2�<��Q~�T}��Mx���H�R��&�QA��zO��i�H� u��]Ru�����(�~����o��;>���^fH.�(�!����i��;+p����;�NUK�ǐ�&�[l�N�N���b�)*� g+�H������J+��5gH�)��jP�z���c���l���<F;�e�E�X���s�ʉ��H]��Y�⟞i�np���%2���J3��<���`�Gu�	1(�')���T���֪x>��ӄB�>���������)�]"|>��q�i��'���P�_��dt�q�}������E�)�����n�t��y��|��H~���(F� _�<;V�MP�Ļb��A̜��\���Q���-�8c��Y≥+t���`��W�����2P1�����瞠c?~�9#%V�!��.樯�1��
�F�����Bʑ` C!�G�Gx3�0��#s�{��J�x�ψ��@��#7��O'5_C���C�X���@�ܤ�ϩ �z� �#�uh�:X	F2�&�"D���$ v=��%�Vيg���E�e�ĄΉ���:P�� �K�F+��P+��=���&�l�c�⟸�6�H��\���c���x���� w2f��Iq�6����jv	w����^70k�s�H6�_���ؤ����$7��]��l@�� �9Ūa�v��~e��?��i��hB��="c�S�hqȤ��WI��*
�?j�f!Z�@�,�=�tg��Hd/&�9��*�Z���E��KP����m��^ќ��bZ�-/�er*�E�ǐO�(~��󒺣���ȑDjht��隱yU�}B/1�J�b��w�]k\z<���6=y?<�6��'[֢S��=tx%���� ��3,J!�h�Q�tLZ�g���#n������!�7����cj�I1h���N�,K���F���C��>\�J,oz;ᅫٱ�<�|�, ���K�E(=�%z>��iS���8M�Q�C{>B�Q&�HH�r��.6Y�hȑ�f��\�jVD����\�O	s��Y��р@�T��A(\ǐܭl���YZ4!�y�Iŵ>�Yb0�����&�� ���;w�L�"t��0R�����?4�x�DR�H�����8D]���e%�eE5|��.՟V�y�Q1 gE�狶ܢ��k���^�t�Yі2�T<g?���9²|��i�ⰝD�N�Oy5�{���8���%���f1Q��m|��1`yb�a��;�
~V�{?0aO�SFj�t���A]�7��J2�ś�f݉O&�k�Ɛ�/�/ Sq�5�QV�1��������)�ϫ��&�u�����-=p�KN\R(ԟ�wH�$�
ɂ� �x`�Ȗy?bQ��������m5�g:b�xm%��U��Z}��}[_�_����e�?���cw�j����UZT"9�Ԥ�?���H�a_�>|��}� ���VZ�`.�=Y;/[�� �u��0(|��u�_����g�����;��|����\ŢX�0��%��>�S���%�Zƍ3@����!0�\~�'���%؀��.��|���5�=F`�O:�(���U�	�ΐg��k��N���LqtZGJ����X�+mh�����Q��Zs(!
�����u�Kl��?9āFu\�]ӺF��J5,B0{�"�R�O��]�q	��ѽ
/����ޡE-2�[I�N%��I�B��4����������|f`���b<��C`�����(Te�W�Κ��6{%�  �I��b��le����v���	�&'���n��-��8$̄[H
��~ł>��G��b��DÐ1[�_K+R@$Hb%�H�I�r�����m]1 $�b�|$���=<�?�*/�#Ji'U�.;���u��9������Z���n��|: w�E����J �)�ab~B['�\T��A<D6)�Ц e��>�^�[��O�u��i�$��g!��j�di�!�pt5W	�޼m����|�i-`���8i��<s/�[��F����x���)P?F�G{�/������)�����N�2j`�E��M7Ϣ'g	�%F"�}�,a�����*�����˺����ܴ
�1�S���p�DS���S�җk�w�C�
�ǗT2��:D�4�,��~�ɔ��ļ�FHB��0�?C��(*�2h�,o�R!�q��Y�H���/�L���]��SM�nP#=L���Km 0Ɵ�b+!I+GNp�޿�Zh�����m �R{�,��eA�է�F閊�c"�o|?(�t|�;T��<7P�F�~
��ts�0�@��sٜp&��B���j�u� h�)�O�Xso�L�ȑ�}���:��0:��k�9�(X�O�v��}(�+��Ѻ�|�1�����{>d����C�� Q�G���u��(R×n'�b�:��il�˜ǀ@�!q��Nt?w��
��S� X��ǽˁ��p5.��*��u/��#��ylAv%M�w	��|����YX��'��ƛ�>p��G���S�.ZH��=�j��E!�V0a"�4p��>K�Q��kc��^����5J�z&@�6�S}<��i�u�NF��"շ�T�W�=%R^����p�)�31Hz"9P0�H���`UdS�^��hta��pM��j>�LʠgD�~�E��0�s��wp�+=FL_9s�O��̚L-��_A�Db0e���H��u,�G��{p�p�;6ߣ�0�/��.�E��6�?���ѪS��q��k�����I�eg�:��-7r�Q1XF���v���F�do�u@��M��dO^@R��^��}�򻷐1GV�=D�?� ����~V�·�� 6�+n�YS� P���7*y �;��ԉ�!�" rO�`ǋwU�0�u�i�_��0u50�,~v���k]{Oh����c,��=qQ�$x�TD1��94T)���`������G�1�8Ñ�K�U��Yv���#T���ub�/���Ύ��ke�������g��sڟ��oN��T�PJk?_.4�e�H���~�a~ `�!<�� I_�*�e0�����{�V�<L�x쳇s��`�g���.KI�O>q�Mp��j��nC 5�z��Ӽ�������W��ZoJX:X�� �M됗��E���WѰr1���6ǒŲ�SC���rF���(�죪v1�~fj
9�sMH�8���ܢ#��R���@�]��7�y�]��Gu*��{��0AOUX��C���z3Z:V�7g�F�HW2���Ӝ�Ty��;��U $N����m¢�c����_{;�s�1�U�'Gp�
ޓP��~���*�C� �����Y���%�� �w]~�km�Opy�v]K[T���Sxy�e.��16Bp8�}g������w���G���c�tV����3xY5J�����J���b�p[- D�� ;%��`�����
������\��'��@	�FC�5	~�l9H$��w�,w�>Ƥ�k�OgXb���5�� ���Q��6&�������/�F�P]Q��FU�I���T��?�K����쯍6i�Hi����j�~cV��\�wt��AgK�[ JE�{Բ%�,������}Q�zY��F���QV���-���C��*��E�	����������2L���כ.^o�(��٣�:��Gք;g	P����y��Pz�:)07_xYeݠ�S�vW�a	(A(w()�6�Ϻ��j�k(�?E)���@�çף�6�%ν��9�J6�9�,X�	N��w���h� 	1kF��zװvQkź�v&����h�����~�!�~�j�Z����|o�I�u*UX�j��Qư��B���zG.ȯ�t��)6����c��ց��4�G�UhH�ʌ����\��1��?�tI6qEvM�Xr9�,U,O�����+�)�H�Tt�t�k�Ě�aȯR�̩��]�Z�p��3�,d��R�0fBa�TÑk��r0
^AU������ʋ���x��ۍ-:B5��
��\��U~�XtU�^���j��yE����<�O�-���ϯ]��O$\s��y�=�qZ.^o�ow�xC�X|?%4#á�12M%�n*��9�M�>���@��ma��:^��U48�e�����CJ��$�������?���Z�`F�̛�^#I��p��җ��xT",��(�L��-���q?�7�����5I�뮴Db�ֵ��_���~��������p����gJ�/�s$[z�D�����ΰ�H��&ӣvX�=��n������ӱè���P���ӑ{�ㆯI��m�H�����@+�25���y�j;A�k����O�s�vJ�]3"7���p`��n��ͤ�{p�}+�M &BJ�1��aX���� �7��:�>Ǘ�ys$f6O[�j
��~�g��Fg�s5)ܿ�~��<��[i[�2=d�����?���_b>�5� �7�C%��]!|���:��k�=t8�I���uw�>�s�{Ƚ�	:�T؛㥻�o��ۯ�$إ��4���JT�ճ�HX
�+�뻈s9Ibnt	�vt��V�0R�|s���r�������ؐl�R��7!A���')��Iun\D{[;����?Q%��Mw���^�B��%��l�z��h�B/�*��Sl7��'��*�j���'��u8{�$�b�ˠ'��d����s�㋝擿�b�����PQ.��+	�F�<0�e=��k	L_��u`�)c�ۋ$����@�>�]W?�}�J����4;�� ��-�?,�qejb����?���1ˠt�oV�,�X���E�$Fiq�#&ƞ�0y�c�gʙ7u�,_+�E�x~I}ح
ugM ��B��Qτ�I��s����m��y�q�� '�8t��#���Ix���`�zZ��R?q��o<�9�JB����6�RϨc��[����E:c��I�1�z�t�/����{�[���E�q(�B!��a`��Av#�D;EW项�M)ЍJyԌ;s��!���Tn��D�DZ�7
��$�t�_��|�	�����]��C�i��N�y㩌����C -�z+
�G������o�r���E��OZ��q�����4�����ƙ�a��Ȟ��uf>�/�M{jkWF\/6���쿫y۫�K��&1���m�T�)V��'P>��B�;cJ`���#�3�B��E��Q���xu[�̔q�'�(ʛK�cR�ȷI�d�<�F�AJ�}������+��o�z#�9ɪP}(�s�F�	���;<.�[��(��=�UT�6�)v*����)[_?4����.��!��^������J|Im�����L�F;^4L�ejA�0%��/�/}o���d�u ����!.m�2�J@;�����:-,'�<A�I�rE��Y�Z�'ִsB!/F7��Q���5��zŏ�Y0:����Ci����������=}h��3�ţP��� 0���Jd��nhd9�+M�(�eF���v��Uo��J�u�N���  ���	�m+�y��XI��m��6�7ayF��:�	H���6~���������4+e��2�Z��X6�E�S��H3P���z].f�U~�.1�R�g��<W��F�0X)�b��*���|������ch��Lq弸E���ч�@55��������M�iz� ��a'�1���1��m�'AA�˹� &����8!(��j�yᢵ�(�5���/��̑�8�#)^9�*T1�d"��9�DR��Iq�R��-�y�P��ЬrQ��ÎE�p��U'�	�	��Xk���&����A�26\��j���yXY}���D���R&��u�S��j8���\����S��Y�6)t+�E`�nY:+�R��"�������^��G��n���i�$-�sh�0���#0�_ ��}z���Ƌ�½���
��6K�=�[�=apQ釵�v�B4bHE1���1���Gk�=+��y�P��A�͖���|K�X� ��m�ZO�V�|��WO՘��MbQxZ)M�Y[Ip`?�_��:4(�j5<\p�
w�c����ahӅ��I�,�:����/*�"��;{U�G��])�wY����9�h�A�=�;/���)��z�6Tw���f�()l�cO��w���k�`�h��?��������XDz��Ν�=�e��%�d�%|�#&� w�Q��s4(�d- r�Rv����d4���/]j�iq��g�����t�;<A$}���r<~o���m',)j�x��s��"ND�ˮ����K�V�s&G�\��̑Ib�l�Պ�J��/�=��B*��𞎛0��X܊8��� ��#>�j$/���8nC8���:��1o&V�U��κ����e�u4�������M�8u�����%������}|{&ͼ��ڵM��f3�� �3"l�b��N^8#
�^x�#�P�(���Ăn��/P�I"����(���U-6�0.H��c%;�GbI>�sP�P�:�$Ig��E��F2_��h��w�@��Vţ�� ��m�����NM��7�KWk�,�{2.�iͶ�T���.9*u��C��A�Om��6���u�~q�:� �ٻfq6�4a*�D(5�5#G��/۽ئ����[t_��eo�Q9�)�U��i'�,����E����X�|�N���"d"�lb��gT6 D0|�V���ߝw�J�F'��C(��/�@��tdO��]�@ہ�D%í�Z3z�ǋ�d�_BCj[\�*�+��t����g��N�����1<3u�^��	��j1-�����~;!�*2��ڂ�����P�nP1�=-���F�43t�m'���IR�jC\kO�介��*�Y�Z�Q��MdAĔO�b�PFt����jwYZ%c*��iNH�烧6	�����F����
���G��?3��%Xu�<�cdg��W�؊�x6������0���|Yh�1�la�=5t����)*n98������P1n
��	�*���h��ݬ�j���V�=���3�"F'��)�[��{���p��ې�bD��jh��տC<F�(��ǱF]y�9����v$�����rg�����)0�:�J7�1k8r��@���p���k��w�������l)wJl�W[O��X1Q�1�1)�j�Ln�5�ӸF�}U d(��l��S�I��K��ˉD��r���%�EnLgf�'���.�H��E�\`��"��3�Ѥ�Ņ�iG��l;�hR��\`z�A��@�ͪ D嫜f~��CmAPD�}�nh������e���Qz�~���Li�������w{�M�3�//��s�K	��Q ���������:��q}�&ud8�gW����	�'k��;�D� W?���+�g�cFc���i��xa'�F���N�L8�7*H!��|�,���q��ۮ��`O�PZ�%#-x��W4X#J���̮�/r.�t�����	x ������%��d]��f��o����A0��/0N���ub����H��x�:V�C�Ilź�����l��n�{$QW2\ߺ��-B�>�"�$&��ݥ/�}������F�3���1����{�:AI羕�{y_;�.� |��?�k�5�H�M���|�H�܌~�.�cR�=ǡ[:TMa���n�8 �[=�F�`����	@[���j1�%���V��墘� ��ϑ��4r�i1����F�y�x�L�3�M5��#̧G����Yv9���`Q%c�����������.V���2p�@^�"��p��=g5D��<�$r�P��y���Z� �b�O��3�̨�^��6��%���7��珑|J��܉���J��#�^��NO��c��i$GR��m~b�-o:}{��4�Vg��b�4w��vz�Xb!�G-���
��w�k4���c�717����#r`��{[��C�)˱!$b������)w�Tȫ�#�m�e6IW|�T��@���_���u���''��7��L�Pذʽ���at�����-�A�/��#�9$��(���M;�s�����?N� V&l���;�C�6�3n�iqQ��I�@t)�X��A�jFj�w�G�����x�uN��
����5{g�e'���ϱ��aP�lmV�=�D6I�Ak�9V6Ǎ�
�3�� t�*a'��t�ȣ���أ�7-I�1VּX~n:}+=�ԌD��X�˰]*�4�=�j�A$����ɨ�s�D6��9��4�^>�̓�&O�c6�r�xZ���Z�`�Kq�!ᘬ
��R�����[��bʁt8'ƹ���p����eζOݵ�������%�� ��HV���������y�_bG�6�\�v��ػ"굢VA����B����M�uѤ���KT{�b��Sdo�uo!�S�k��E�80�۠I��G��	���O�<�*�)��7َ8�5 �,�,�u<�������D�����r!��e����)n4��e'����#��+��S�rG~j�J��6V5)j�E�����c�$bLyk���vX��Q��Ď�ωǴd��lS��)j��_�\�$��?�i�9ì�_)mG�d�9�m�ӈ	�r�5�|a81mh����!	���tfS�h��R�:���r�5V韟?��F�^b�2+����ww����]�*�U���sR�8��$`u��1��^m�Wv
��4>Ť1�;�Ɔ5�џf��yZCD5�-����Η��BWV+	f��*��Y͊MH}�.qr���S���Wɇ���j���7W���-*F1,�w��M"�����Ha]��{o�`Zp�%��
-�DR-^3������5�,Β�_�4�+^W��>�c���G=DJ<�$�|~�u��]h��*�词���i�:`KaCC�����z�������f}�\Un$>�{�ҿ�P/�tR�9�>�V�h��T����i$�h��{����{8�0�ۄ:��x�9�%�`���UX��)����߮(�@�?1����Z��J��h���:C�R�� �>����l:8Ȧ��4���J�L*	�]^�]'�����'����6���T`�I�Yۊ��p�4��;���uй�y@ajc[���U1�\��g
ɯ}yɺ�����T�q�<&�l��}%�CB����~��(�]c�˺UZ������	oW!v^<I��Ԥ��w3��#�S�sa��`OT"r�3���ǀ���'~F��k�۩'i�U�Q���`׵��,�Jj��w`56�P�FVCsD�jʔ�!/�ȥ���`�	�-m+<(�x�,�����L-a2*Ѧ;����x�ZD���u�y|���`��Q�w��Y���]yk˿�#b�"�0gZ
[xT�Y�+F�t6���%�Y��T�ήa�^|��B��s����Fr=��PFvͺz�����E	�x������/��f�?[~}ph�D�T��d�?����ڄ�~]���������K�a��Bظc<$���B̻9�륋�yEخj�"���u�)uy�ޥ>�na�'}�W 陫�y3��m���
G����� ٭�a��~�9�L�C�h���'Ef>7}�R�[+H�҂?u�3;O�ϟ y$� .1*M 7_��s��ڏ���3�.9�
Q�m�i%���2����e�\
$���t� HQ�!�ʅ{MՒ$������X�H�>�>gA"���d�?7c� F@6q�'�m�C�f=�8�6�������$O�|�rw>h\����l��Oî����VL����E�)g]�����p~ՠy�1Ve������Y��ǃ��Az<?�p>!?6�	@�C=�,R��ٌFA��p��u����Z7C�:.&������)j�K�*����Bk�NՌ�.�"���(k.p���b3,r�լ��@�		��;��XU�$ԍ]Tg��`�$���n$� �3]���^u��
��o�aL`�UIgl���[�ɇ�`�>���5F=�0,'���V�t5�7�kdX�����Q��I5B���slT���A�@C;#�РRY<3�=�c��}�a1�2i��I܁]�sǋ��Ym'U�8�^#�'�D�}�S�I��n�ͤ�_(n��'w��"�����	*�F���r����.��eؗ. �Sa�s��hb�6�>];$/$/�5)<H.�V��ZGk��;��=����8;ev������X.n�dm�9~�%lmM�I�}�A^��a{�f2V��(b���Mj<b�@��2��S�q̘�T�i1$vW������P�C�ּ��&eͨ ��XD�(c��w1L����y��~8]���70c��| �5�
�እ�a��7��0.��i�XUpҪ	�F�sO�� �*K�}�#�xtW4�VWF{�㔺�n)��n �U��q��-���-�'�Q]����ā\1��:?`����f�U(�t����օC���N���X.�.���}|��>�i|3�"0��]�U��`Q9�)ýP��zKr�m�I�C�m�A��v���g�*/��r��f��I:��WM�f�zK\��5�i�N��o���� ����ªL 0�����'��ja0K�y�#��I�����'+�ҬR�EO�A��c��� �����f ���椘B�إ�N��Wiq�֒:oUY��t����Zj�]xM��1_���Y�G){�3������
R%�S�b�o%�7�T I��u{@�44��Ղ�ߌ�^�P�`UǺ�-�J����<��=T;�D���k=5R��3R��dX�L.��T��s�Q��y}��M��J*ys�W֚��(9ܺ�y�� ~U1��҄-;�;��~�ӡ]�'������� �'[o�5A&Ae�"��`���KN��T٣y�9V�;r>p�>�)�/�o�e����z�Փ��XC@pq��V�6s�e���@�珳:W�=��_M]$L�Z�!ي��5A��T�A-�*n���*%�#�u��o���ċqbK����c.��L�K�H(��rkg��kԪ���h��N��n����b��O�̍;�¥��`$.������23��i����ˌ�����R��h@����NJ�5���"G�m6�W���s��� f^�Ԭض��e7I*��_�$a�IM����K:pJ6J-5Gt����]��:�'��z�ƨ�;�]��j�9,���t �oh.CBiC���PC�i:t�+] �2'Ĕ9mA	~'XP�aMΩ�� �Wz;Л�Le�{����`ڼ�]�WpoJ��G�3�E�;���˝jo�=��7)j��z�}t�i+��7�'aqG؏��-���{,ǎ�x�U�^�6���9B1�ܾ�h��;���ɾ?n�&n���c�.��Yk^�6���Q�X��E�.�)"�
�����f �[�ɔ�Cl����_'�9�����
Z@f�(�������G�:o$������wGhԧ[�B2�J�=������៦���z��s����T�����"��O=�X.5��� �`5!7�.�u`���J�ea%%�B���[��£����!P���5�׊p٩�B�{�#Ya��Q!��a6�p��E��yQ� ާ�ϲ�K��W�BoPUˌ�"�Y��e�z��Bt�I:F�,��hV�����kl 
co�[`�_A��n��b�݊�.��Z(�u#���D�=��˟�M�E����^�佽*d7(v�e��y���;��bC��B�
�bĮ�k�Qԡr��u܎����8�|�N�1��0T���61���>�
��5���@$����ı�=6��U�{=��H�GBVw�|��ˎd����n��S�C�� �Ĭq2� ^#���N&��go���yP���v�!�%ƿ�;������r��f��(��آ�k\��AL���x�GQr{7��2��:;�?�Ƀ�S~��������Y ��Z?{|�
�2������y4!FS��p�ݯ��`Oi�aDI�YLY��{�l�"�@6�p_�d������C��B�:S��Ϣ����"�[��ʔ������E�p$J�+��'�p�]!�� Α�Z�,�'�!4�ӷJZo���a�}I�׷��} ^tQc,S������Zu	�M��Ԭe�_�ˮ����|�=K$1"��H���n�d�4-�(Î�r�J�3&�Qh���k���J�T{����$#��k�+k����x;�]��[(���qIbf:���	熈 oy��
�ez_�XD�7\�w����`M	\[+Y(T�Ż�`X2�-hr�v����1h5O��KԬ�ږd���kO�����%�!laHV�,V��b�X����шWWl�����_�5��ճfg��+��Bˊ����Zm���nS��k`a?YBm�K5�o�B�%�/�&z���j�*����2�+`���:�&��|��!ig)��%���.]��/I���	��� �e��X��H�Eț����5E4�z�%�3T�e��I�X�j1c2²�?y�yq��I
�ϧe� B�G��u	5��h���>��}��v�J��HEŜ��^^]��Z]◼v�O�b�
�:���	�������:~����V0����
��y*9!ٶ��9�&h�u���Gd�M��{{�*��Vm�c<{� e޿M��\���AK�P_������X�X�̽��t'M+�{��;^]M.��PT��!h���q96AGm`i�R��(6�;�zk���,D�aw���74�z�/$���j?�Yl8]�� �K��~�y�I����w]�!�5\ޢY�8�5Y����Xb��Op�~OO.U�O���a�Z˝�5���zp~�[��[ ���s����C�,u�TZ�F�[�q��DZm���	�ͪ��3��o#���z���m�,�#nP���UL|��Y��q��a�����熵��ۉ�no���B���۪���3���������h�R��*�ü�M[->��s�։�1�%�@n#����+�)���+���<��Tf�d&q�׾U��9\��#�݅(e�zuI�#$@ж���.��#2�a�H�����Oc#=z��^>31"Yk��O�ùþrѹeA�RrO)�#_�W�g*Dr<��M\N9Y�@�UT�A�`^�2 ��~1b��	�-�8��b��W&C)>n�\���P�Ӱ�Ȥ��&Di�n�2YIM�f�D.�l��~�oG�ȇ~K]މ@���,��=�E�5*��IK�04��ٛT4F?��c8���ӧ2��ΏNvfB"3�՛z�a�T�Ԕ������a���s����GmWdk��?2%�\
(�������sI�ET�Rd^nO|(}j��Ўk��E�'���躻��'�yL�:�2W�V?�6�aL�qX˫<�O�y��8�ꡉ�R�R��: ��!�ᗚ��=�������j��θtzT���Qk��Ro�|�C���V��\F�!rdg˒�F�&��8e��3I����U�b��4m�"��� ��n�޲u��V)<b(=�%9	��y&�����@���Q\����8�F��0\�rW���=��tɻpt�)�)�G5S��� )�����N�wi�	�u?�m��2_�S $C>}�uayU忶	�\{E66_�609Շ��y�j�h짣��)�=��7���oכ�&i����N��l�ZD��v+��%����Ls�r�a{�ǂk�����5�eĤ�(�8��Ѝ	�C6�3��W��@�}R���
�M..������tT��X	���&����cz����e�'����8htď�Ѩ����و����g���Fv�P`*׷QFI�q����8�w�_���:-�P�1���Y
�SG"a�O����`��A6�]G�ޜ�%�3�kb0�#ԏ��%2TS��!o��/���OA�l$�c$���� ;�ʄ�˶Q�(�%�|�'r!ôa0���6��T���؀d7nv�+�۷[b����5)8�믿�7�.�+hW��n��^��K6��*���`�E噺0x�К�Ym����ꈐ��7��T���J�i2�Ń�q�?&�q�T}��jt�(�5����wvV���������6NIJ K4i�{�e�J9=�c���|F�P{kS"	4���U�X�L�R��B�����Q��Q��j��	�����\�8WS��]�$�N�dWvB��_咬���ٵ	���/$m�6��0]�P����I)o��W��?5�{�8�xͬ(���P�V���-�n$��<����Ox�B�֨�>�*X�,��-n\�h�\6�(��.j�H[��_�Y�M��ܚd:\��?�[R��j�����b��g���ǹm֨�D%a
銽�8�{�>l�G����U}�Mmmf��	]Ζ[�)�f��#����/�ii��a�'�D�!������ja�'����"ؤ�{/�+�0kyE`i@9�3����b(~Vh�G�CCtҵ5۹��M�쳭gP�n�����	��$�݋�ڑ�d�#,6�c"Z�Y�N�1q�}�iLx�K؆�`n�����pH��}@b̚+k��毭��ŚCB��ٜG�Q4Nٵz�g׶;�h�ه��ӡ���Te�n��i�����k�]�"c��}>3�:@0� ��P $h1܏;0�O|�Q=i�e����p��wZ��C%�.y��^��x�Y��L��e�"U�Fh\MTۀ�!G!�
�%S␥	!g�ࠟ��R��G�����)�!8eb�f;u�.�,\�l3?����a�ڙ'�~Gh�-����K��15y\&)�%��Jg��AW������#��7i���NT��z/R깨�O�G�[-�^�*�U��? ���k��aĐ���s�b��k�N����Ă�(�}���!MB)`�=�8]���L��LÇ�H�$�E��ř?`��U���oo^�1�9��Ů�����7UX&�� ��I5ߛ�6�%����w#|@�e�ߏj���eDS]��ԖG#�dvj\c��4uMH�8���L�O�7ڣ�zG��v���v9R�k�~��Ǽ?m��u��," �����3�L�$Y�+���+~�
��'su��w�.k�
W�����E��)S�w�i����hNs�8j���,���(G�����F(#/%��d�@�ڽ_�+V!�,�M9��	0�����JDob� �Eș�+YQ�_�|vm�o��2���iw�u���)��w'��vc������)[ڈ����~��5��[��zU����}�@��d�9&o��F6q��6�W�;�}�&}S��٣�i㗨��s���o������p������v�5"H��,�ɵ�&�m���dgG��1f�U�Bdx\7N�����+i����:H⑔y��;�r���t�f�_ E���y�h��-[N��|�]��B�_�Y��ϱ�(���]%��D�P�q]�8e�	��?��=FTV�
��Ǿ�"s��wU�-܄�@�ڎs�\C|Ԥ¶gm�1�ϰ�A��8�K��`P QR��vTk���ZN
ʜ8i�s5+��Е�>��V\�7�pH�_��������Ye� ��[ʶ�׮��mJ-�������1���_1�5K ��������e�H-J��rg��xtY-^��~�W7����`|4��5�)����H�����	{����=��m&9	�'�f� �l�`�����\v@4��/JO��������+��e>���T=ग़\�v���I�IwkBX��7�t�(��s�
���iT�CrX�ݦ��وp8U^6��k7�ĢU��!��U�2y��zE���m�Q�i�!LC�A�����RN�&�e����=z����ƷY)j�r�������H<M�A��GKZ�Ϟ��^��I�H��[u�l���f.��\����CGBV�ck�Gmia6�^k��Z�|�i���8p�F�׵U1�N�k=�f�3x�9O6��%�}.��ʔH��8�m�x��3�5�ך��Xe�@J}5=!�(	RR��J�c�!,5��szT(O ��o�4f|�����K�A�{�q�g�l�N#.�Ϗ g���cq�(]�]唳�|Y���=��:$|��JH�RO��|+�Ğ����1yߢ�����Me��o��@�e�w��#3��&��;��Ua�m��-H�U�vi��1�l�T�����R�yt������:�Il��Zjⶺ�e{�\0:��f�7~E�-L@S�gsv���'c)?_"��� �aZ��W�}*	W{sEU��R����5v#��/�Ա��hD�%ь�Q���O�c��@��V1��]ސ����]�qKp=�#(:o`�l���z�GH�r�X�ڇԌ���?�s�X��(z�]yB�-U��&O
~\�b��Ɨ�a��PJ��M��e�:���z�⥥��&c�k�T.7i�����5�P��ЦUO��˷���|�i��>8T��h�s��$:�N�5��9��>�aa�6 �F� ����abb�E�O��?��M��_@}�s�ؓ�
RY�#7�Y���MG��@������y�j9C��vr���Jn蝔��|����Wso��P��U��
� �wyčV!����4k_4v�1�zB҄z�NWj yFX4n��̍y�j�[V �¤������٣�!��Umw��V��?�{�&Z#I3AFHj�,C7kC�V�𙏅]�����K�q�^[�D\.�
x���`�/$�\I�.Z�Z�q�Dp����ӹ�r�[�J��%1�ܽ�AR������7�����GC����x�+'�����{F��B���J:j^Y�:&�(�A��̾�������$�<�J�.�+�ON�4o��HJ�)a�_�dBs�8�������	X�X����׎mr]цN$>ų����Dw8Es@�o��}aN�~6Zc4*D�qww4�j�d����o�	MJ�0k�����(���xq��S0����ݹ��i�k@b�%t���:�zs�hC�f�$����W�����2�&v�s�v�Gi+�QQ���+�NqD��e��JV!�l��(��A��!�6��6G��1a��v)�H�e�F�VZUL乭��昃Zlv�(����?��=P[r2A���<��FG�i2����~��&�w|x6kZ��u@�xqȨY8pp��R5Y�AӁ���JЀ��6GGк�7"��"!d�-�ۀN\�w���pVl�VP�5��;�����Q���b���'��2)Lfp��)o4QAv�����_ޜ�b56U1�}��DY�L]Vg����X�����gN�>��>�'+�F� ��>�@<����ཡ�1�֠�]ק�.)�ˇ�DGc�,�>O��^`�<�N�tB���9M[�`��}���������g���nֲѹK�N��$�1�|!('�$;�ZKq��X��	g3H�!�!��ͺ��ٟ��\	�C�lۍQ�&o�g�s��>_ߑ�zC#IR������>�n��<`֐¢24�U��D�A��Q���<�[+��~�J���RX�0*��7d���l?��A�@��v����=+Ӎ���Ү@�ݕ3b�Ms�e�A�tU"KC餑r����&#�Bf�n�f����/l�=�����3�I�,�}'	��7�����C$�N��)g|�sY��	(��]c�@���3����ޓ��2A�,���-��V� ��xi����3ل�h�$� ]<� �>m��9WrX����޸?��O�HEI =�	���k0���4,#�~u�H�\�����n>���,����Ix�:�:�nх3�ڐo���+2�:���䱹�.h��i��:�j�:��?��ڏ#%�+c�8��u��?���1�ineϔo�3��ׁa���"r������D�kL�W<�KC������>6R|/IiL#�hk���|��S$֡�h���n;���x�����q�XmV�f'��������4%GMK:�=?����wU�l�'G�KhNe�w�8h8�l�)��q ~��I9��{6`�_3�����/`�	A��M$�EdB�Y�2���L�٧/�X��|@VN	�p4a�iЄ����x)�'�W,1/l���,	�N[���wT�[r5�,��? ݞ�04��^>c�'+�c�����(���n(���E���L��C�q��T���=#f�`�.�����P��%9���{!Ö[�rB�¾��
��Ԡ���39����F�����k�!�yl��7 �Ee�g��bOC�xv�o�N�ƭ''��Yc�?0��) f}�'=�N�p.��RJL���[Cj�E6�YN&�_K7%�B��\�GCSD#��q�����؍Z`�7������*�ɤ`���}NP$�|+��s��"/,�%m�I�P�u�a�~1�O2 J��,h�����Y�1�����q�7KJ9tz�G�]z��*6��>ו�|���
�����z:�s
+i�,�%�������7�넒7����y��$�u��9�T�.W��ޙ"��6�;������rS�~��B�H_##��&w��)�qo�p�Ie�������]��pN �$+?]C�0��֦���]Zu���β��9���7����4.�С��\I<M�	�9v����҇�L��g�>������Ҭb�LfjdZ����с��Vx3k]�/&U������� K@�/�8�4���mQ�O��띻����� ,�2Z��Pę��d�)c-
�z�-7c��H=���{��F���MW�?y-�K��L�%�˱��0Tu��=&ݿ!Ks:�*By��k;�����?g�3/wh 8�'}����H�ξ?�
G�|6z�v�^�åB�D����N��?����&dɒB�����ߋ���	�_pҭ������;:U"��:�T�۞�'<Ϋ�ܢ���l�,j�#ih1y�:�u�ݖ�teٳ>��Ƭi����bS�<���I	�� ᦫ�<^�#6��_N筴���TJ�c���������\�G�0�'J����`?�+�]�7~�iX��,u���`q���A�R�fۻv7�BJ� dkq&B�+�}���W�,dtqZyN(��Y&���Q.��r{�׌\f2\3d�T�^����-��1�'b�[�`ޒ�$'�����ISPXO�2�V�9�����r'-"��!�xM�+�-L��լ�im~w��9�,�½�g��:�h*�4��	�����q��y�FmJgwnB�C�54P�+N`�-�{���di�T_*I�Tͦչ��s��Z��UDe�I�6op_}ۡ)��i��Wnus[B�v.���h�s$��0�Tj �����@�zE��yJ�C�*�(�t*�����Y�{�0vY�L�}�=�M����jv�*�V����b�{�,��V.R��K*��{I���G����UG�i�� T�)x��+q��^�?7�'�ՏY�݆�U��C+���Y���x����^B1���h�@{`}�Nϕ�Dg$ψh����t>�PVխ:�t�ɇ������R ��F��D;��#���+��I=�K�Z�q����gĹ�bc�lb�P��8k}t`Ia�{E`Ɖ��Se*�^U�<�%�+>jX��Q?}R)��L/s����؎LH�ϞfΧ�إ�%�f�����`6�'e:��9J��1�g����5��p��_)���E�U��@�vPM�S��{]u�%����_Թ��]/���Q��[�m�N��ۇ'�����4Qw~}/��]�J	����j
��Z��t�5~?�{�|;|�A�Ϡk���)57�{���Ҟ=��oi[b�k�7"��k�L�ڨ���7��I��M�6�F ���	NL��|o���٨ʗ�<FD�T%�dϬ���s�e�����G2�w�Oy<��J�+�2�=�[>��+�6��9��P�)dG�,ʢr#:�bI��F���}�i0G� O�	�Ά�S.-���,���Y]�+�8�<8<5j�w��,�Z�ћ�J�.zϝ�1����2�i���U��$����K�A0�?9ȼ�?��^*q�. _���)�V��VK/t����8����\���K�*:'j��1���(.��m�vU�|&eD�g3�z��H�6��!�Q�/
�.��E��_��ȣE浄��[Sɨl����w	s������?ۇ�����Z��1��W�BB,������V��^
~�P�����%\kn�*̶��dzr"�y;�NG�,�1|��!��=_���iRR�+�0�`�bBv#�!�f�Z�_w-z���A�B4u%WÜ]����A7�d|g�>��M�zm����xÄU���:
7�����9F�;�j�c�ۨ�ݿU8��xވ;+��m Ț���a��J�t�}�Dz�T��WĄ�P�Y�St ���'b=�zTF'x�ab�56��f$��c�>�&�ry�aߜ��)��z��\B�xe<4o�ۿ�gM��W���4����e�&C7��}��DԊ9{��E�$h6�m3ly�&ʑM&�b����v�f��VS�����r K5f���`Y����AR�t�/?�Mΐ,9�tC��"8< ��8��y�+iE��x�0R	e��!� �4�vx-[��M��G���U�05ɲֽ���~_���|-y��9���(Z�D����,/¡�=c�<g=jJ�H�lo�w���;G�����k��S�E� <���6�a�!����bo��}�I�*��mKK�R���1�>Lp�a���p��o��$����(Nɡx��=�,�%����;,�t��1�ܸkCG����9�P�����#O��0�0@���a��/����y�C�Lt�N8:�<Ȃ-�E^����,]Uhx�\������"8
����gI��S�P0'C�Z#�D���M2��Q���<�2m���B	`|�l���Hʂ����EY'���Kl�u�|��;f�P۳rƣ��%?����6��<�P��s��O͇��.�En}��&D��s�Q�������i{]�\#q��6�F1�����4L;�-��4k3�#�Wf�W���|&���~F����t�i�l�ޚ�	�.L=Y+s`�c�j=� �Ϛ\L���|-d�a�r�G���{՞��b~���Јͯҫl��d3{^��;��tK�+ ��iV�gV����5�e����r@��^�Å��
�~��ηDE��Rأ�{"_��@
.k�����!}���)�����i�w�c;F�����&��W4�|s��
��ys���Z劌of���[�I��ߝ�n�&�a�����-1���?H�|�7�F�7I�7
P觻�/4��[
��3�#c�6�syu���^1��lR?��i���5��Gmy�]ut�[���E7����O��-�K|��<���]+�$�&.�K�,UHSۓ��q����ߝ���w4d�ad����'&�/o�Th,^}��I{�[�W�K��b��`���P&�~nOVjZ�z���*��͌��bL��[j5&�ӋK�K)6!���\'9R���q��ZS�}�rwJ�5�̻�.uR�^����F��5"$Hh<��dWQ�/��C��K�ⷽ��6�
�C@+����'>��Wp!k~8d���$���H��N&��3@΢ ��^�/C�ꌻrFZA���>��4���Fo�M����og��~����B'�9�9���W���K�X��J���ERp?c��M��}�ۍi �HP�����l(�IM���s�1�f�EZ���җ�lw�����/h9m�aU�T������C�Cc-܌K�;a^[z�2Z�H�k�Q�m�k��A�>� ��E`����w�\G��ͣ�/ۄ��ܭ��i^Is��b�R�y ����6�
�5�f�2� .�B�ό�0�A�aq:���=-��-�<�O�P��d{��
7c��l�އI��mCR�����{
d�o9�XfW�4<�QO��¯%W���`*w�B;'m3�Y�"M��y��8mK��11yX�zQ5��=ȇȼ���#(�tLuެ�f�ű�<'|�Q�i��O�6���m|CeI#�����4�lCZc �[��|م�{�%��j��m2	�� ~R	�d*�l\ynm��_vWo��[cA���>�W:	�9B[ o���W�������x�ƃ\����9��=�.�d�@���>~FKB`�F�S^.��D�T���2D$�s�����+ų�1�m �)N��T�{���jUXx�7�B5ϑg9+�L<Z��!��$b�fu+�}T��*q#������-vW�hv��e�o��/I*�:�a�;��z����S4>dU&<>_�P���kn��ET2����&�8�4iێ�+����=�s��$.�C�ƻ��4���f��P�4�����2����[��ӗol4M��3"w��Is�&n��$«A�k*�Yՙ�%�|*�s٨�6R�v����l.�AaЧ �lB�^*j���ꬁ��8�m�����JȖ��5�UY�!��П<,:����u����Yu�=�l;���0~`�C��>����Pz�;�2��T�v��]`Jh���@���o�l���ɜjr��d�K�	s�Ć�[w��)�.[B{ᾘ� ЉZuP�b2>����r����J��ni�!Q�PRY����GIG�|���v���c�S���r�vÞ���p)@�Q"O@F�~:�pV� 
@河�r��ӥK>KΒJ������Ep�_��}ktw�/sRs0 wj�� Z�-b* -^hT�[��=���~0E��q�+PB��S1�q����˾M�S�gUN���G+�h�{>��Hg6�]�N� ���!+���[��S����Ҹ��ZL���(��e,�<��,��Ȏ�$��J	�(�g��#z�1�ut� �^�}^�MK�����CHnv3ka�[�,��;�kb�a80EZ�^!:d�TE��t_��)8�ն@��ϗ`S6�ߍ:/-�hX7!8��mOK�~��q�F��&�!м�з���[���G��&.<��v}­b�?���
��txw�=�GK�,%o�{��Z}�ŮiaE�q&�+��}�5��/o@3i�S��b����j�m�7jr�-�ׇ��DS>K��Z��'��L������,˛��P��ǿ��[/ǉ�ǲ�_y�ά���9d�,����4�1���<�&�����o�R� ��O�2F��.�}�9�,��l�0����|!�q	:����Ĵ����W��ݔ^�����g��{=(��H�XXS�y&�2ւt���j�\(�s4��Ɣ���-Ӣ�6�>�	�U�q��7u� `ٍ�Z�&6{`�% ���`�A<�m����<�{��OHbD�^��.!Ν��[�������������MЏcXކ��n����?�����+�S�=!��ѣ\�u��7���o�{i_.ʜ&{�X+���S��,��[ۃ�5�1��
� &K�ߠ�,�N:/��ެ��Ѯ��Y4�J��fz迨,�N����c�4����w���2`�⟆�
$�w�kD���0���V��74u+zB}�e���?ϵO�"~�ok�7FS�Np�f����2w�����g]7���s��4�3�lv��ȓ��ʗ������dI���rɑa! "_�X�C��<�&�g�,���$�u^qc������fx꽏�}������I�h
��dv�� [C��Qv���a?������i�f���>���4��_ڀt�'̺ l-���"�1�n	.̱U�`��4R�p*]s?\�T%*�R�c\H��?�a�nS�Y�ȋZ{_h)0&��<wT�M�M�r�)2R	��2e�������W�x�k�9��M����ݽ��A�,�,�0��ƿ������-6�DCR;
H�&�<�[%���R��yM5�W$e�2����S\�h]��5�)�m
û�p22��
C���o!x�]��Y��?M�,i��3�"Q���_bN~������N0P� �Z��UeoWgF�
�`Y�-�V���19�Ú
 T􌈃�%g��/�S\�Y!�@=C����������k�B[X^Aڤ��GM}�i$�M�Ű�d�����X����3��鲄��zO}�?��Lk�֥�.jU
�>bY��_6T`ʬ3�e��}�e~�� ��b9�H�C�x[l��)��+t���� ����=�������LZ�F��	)��Td�u��VBK�k%z�z�k�o9-����[J��fr�^ɇ�,�0Mi�ay���C�my�A6�|
YEN�<ϒ��C"H�B��=�~Iu"�H6��{��0�P?5�s+��l$a��͙<���x6�7�}�hפ�4����!�����Z�D�:��ˋ����4ȯ
�N%�����>5U������h��Vyi�kW,;���VS��5.���~��	Bc\�	N�"�}�UTM�p<��àpّ�
=�h���	S�E^!B��s*B�{p%����.��0�����w����U��d�4T;ԝ�7&�����;4����=NS�����?rcBw�]v�X�5si�Ƌō �0��+�e �$[Dض�|Y{�辂Т�9��UD.t�G4EK��_�W|Q~P�]�Џ��^���(@���d��wp���_I��r'��O.ФM�%�X���خ�+�4\	 tCm)(I����س��-i���@E�n������I&��%�: ���Fr��A]���sQ����`&U\V)�wй�z�hΩa�w���{B��U�zJ�Im������[n����w�2c=�ա�� 
#�n�����MR^2�Ж�3w��+Ѝ���m�;��Ž�W&p�8j���2Sg�zRR2�@/�7#�A~�!FbkllkS�����
_Ո㟩:c﷾�8AGr'�Kċ���@��ǟXWX!=c1'�ݨ^�0�Z[ �E8J��2"{&B��	�n�.�N���OZ�ǩ�5����g&$Ox������I���ek�J:�A� ��,=#SKmz�K������C��m�b�s��v2���u���F��H����"D��@�ܝK�ư	6aOe�{l�]�	�-e�PZUG��q5[ ���1<T��/��hq�{�H�댛g�1�f��듆�Y\�Pa��P��}��c�� [�ۂ�3*��S�@f�?�r�]q~�5ay2���2�i���4����UI�h��7�d��MxR^;��(�R��Dzb��[�~���E:��d��z鸞�W�j�<�xVh���+X�eN�0">?��B1��D�U�ì�x���i�'���T���k�]�1�@\"���>G�su����/��Ha��F��ҿ���#�G�9D{�R�y#s:L�?��3�U�O.S����4ʑwa^�J�'��	�au�wۃ��A� 0���T��\�}o�m�Q4��:y)������ǻ�F,𖿜�kh���@�K�,x���L�Y�I�9�Ѥ��K�im ?d�ܫ�eu�����%�@"� �B��6C�PN�A����e3���1�C�Oٽtq���\[�����܏��!��KY"p�1rvk"C)}[��r?�ug�����K�.G��yO$�4e�-�_'5��Vj��¬�s���??��ݏ-�Ȏ��5_,+�~�����9�UK����?Q�B����}�t��Q|��c!�Q8F���6u��ji��h]�]b^(80�N��(�^��l	ve����8�od0�,C��ig5��(o���������D$�� �I �^m�$�e�]�v�Ǎ*/9D�_��?��P�����!3٬�[a�.�X\RlĚ�2N�Zl;'2S�>|����;���aح�}�g㝓 >k�x0N���|U_�٢��3xk_`��x�|3��k���j`⥶�Ǘ��$�'�:�{��m�KjyBu�'�6���*���^(e�P��K�ٽ����z(q�C4��תL��a�_���7c9��焀�1����-��P �%�?cI�?�m��^���WP���(S"]H��{m֝�su��"-�]['+�y'�T�8-�_��b���wnQ���:P�?��`1O����B횛���f�U�?,s��?�&#)�S�j��^�+�"�V���pӍ���%߻̔&4�����a��)y~+�I�w��r*���c����C�E}=~s�Z9ۀ���uB�2��D�x���N��eڦ���;ʲH��� �Jd{9�:Ǯ��Ɏ��W�~?Wf��2��`�J�e�\�jR��b�݆������~���}��5W�����#�6"K:�EVl��l��̴�Ef_ �+�J��� ���g..v(�>kF�lӷ{i�MO�I����v��{{��y����8V��B(X��Z��̃g�����c��ۭ�ݟ!��$����"�]���g`�:�O�ȩEθaLlYM���s��;�X׫�g�Q b���O� ���"�����+�N�ʔ�8�����߶կ��1�@C�M�*T��}ݭW��ݾ}�yH��}�q"\�U�ׇ��6r�-�Ǒ��L�S�B]MZN�)Q�!�|�Ojh0U"������<:=^7�P݈+Y��ޏY�'�/κ$m�]͔�Y���2�� ���'k"6���t�� ����t���w��J�"�s*-\�^�h�R�1	������ ��߷�S�`��ޒ�HhM�d|�g֥lXۏ��DR7Sqv��B��D���V~�T?f���J����k��i�-:w���%9��&U^_aV�i�ɍ���IvpQ6�% Y�J���Fv��8����]�E���Nݶ��]���D�g�O�Pҍ{�
C.S��*,��K�W�#p��iYǟk�'H��!���9�+����-�pz���G<r\�R�(7?
b_Th=����ع4� xS�#�@=cZ��r�_�i�@�A�Ɓo��Ϊe`1቎�q=��l~60^̭���3M7�5�O�ޱ�Q~�����x��(B�+W�%-U����u;�Vծ &֒��o��J�d��{�N���\X�����S૸:ſS	m��u�ֵo����܉֧���y����g*8�HmSp��9l��d�4v�,N;�'�v*�W���d��m˺�7� ��Č��E����B`v���ă�Wa�DJzIw�Ao�p~��-�"������>5�5��_&�W]��"�a�� �]�ן�.A&�@X�1ǚ���,�O�:y8$�!���]�Wq5ɺ��_ji�!belH�NC���p���X���mX~�3B	�=����+i��1v��Ν��~�3R�����#�N���2'�ּnE������ks4�����,d�Nx��.=��*�B��&[�69W�Nx[3�=���N�Θ��m)���ꠃ<��Ў����ۥ�JpOj���pF�
m�{0T����=1i�PJ�����4��O�-O�"��Fݖ��u�%�Cg�P+7��Mz�N{��F��N���� .p*��\wΌH~S`�jC��C�Ǝ���ĕ鲎�T�o�&Z�t��"�ء]�� ˮ���}���Ο�!m�@�`�ؽBZ�ω���?s���j��t$��	y��	���rI��7�ا�.lu��8�:�<$�4�T�3V���G��ET�4s4ߙ́u��Y�U��R	�NI�*:W��[(r�4�#���ˇ��p_����_Z.${��<�����$�_���9|�k�'݁�Ac� ~��AwB�=�Yؖ(��Z�7f�>Q����C �J:.�V�u^W�۝��[9�\�UN���#��%��\��,���܇�֊����́00��  �����Jw��K9��Sm`J�d�%Ӕ��uȹ��`�]h�Ȼ=Wd=�᫆�mVC��Lͤ��~
��n�/�{��1�Jm�I:�1����'}���c��^��j�s�S��9���?�0�
�k�.�Д{�nI���0�Hķ_��"왇==�D�� ����/��V�xG�yCj?�fiR��q�b��Io�Ml��k8g~,���B<f����*�
�����#rp=��$�R������KΓ���Y��䲯%�J��Y�o�οOc�� �`�=^O83�|&���4��M��ؘ�	W����S]��
����DR���$9 )Y*UF����-��"�����4�-��b�c�����)���cF�1�~vt:�'S;�+,iꎗZ���^$j h���<�$��^IS�+|�v@����;VR}"�bK�J+�� \d�$� �:j�Yd�xO�k������h�*F�W�ѿ)�Q�	=&S}V�^��V�>!�����
�Ö��[��|��V�2�"�z�Ð7�N�q/�	�������C�����&�K c��?M�������o׊˕0[z�;]JGo��d�5�������i�h�J�IG�ǘ7C�ዅ��$���'C�r�c��hz��1�9�����ˋ�x+��s%�uo�U�h�뼕���І���Wռ����B-m��3X�2e4��
��Ի�^����Z�������Cw��9(��@{
!�θwOe��0�r���<�=�=��k�b��#��	/	�,W@|���6;b���?�dmωG���|��EM�pc�{� ��::��ķ�ś?,:1�����-p���V���dRǠ�����Բp�EY�gր`�r����$}yV�ѣ�ĩ� p�C&��Xf��Rs�����˼cl!U_�W=�?��I���3X�%@������
�(Ɖ��V��]�Ԇ�h��R�1-�:s��U�
�m�3\?ӳh��u.��A�5<�U_�)�Bi����§ 6��ͱ榴UV!-B�T��
�Cm�����O����I�T�+�2�!4c6Z�����&H.���Z�P��;jC����W`���'l�yፒq�Tjӹol�{���&M	ؿ�V��YoR0���)�(&+-���؂�y�2��X�P�Z�S�����Q����ew8`|�j����;���XF ,��2�����u�_XDW�>�D�h%'���������@D��� ���4ʿ;�4D&{��T4s�]�9�d
��c��
J1^DyRs
Io���g�ޙğ>PϬ�ck��,���G*1Y*��1;�-B i���� ���=j�c���"����%�j�zsG+u�h�:�� �w�[��=�v�{��im���xl.�Fϰ'n����Im8���~��Hg�
;�#u���C �`p�Z:^]���]6���z����y�{h~��s���
co���oܴ���8ly����Qw�wt�)`~�����KM��7R�"��鴝f^�g�=���`�3�ۧ�I�<�Flr�������B��ϝ���c+:�h��:L��W�N��r*�rO�br�͌�����1�\\���Z�E[	Tv-{�oLGԭ|���t#)��fqa��Qj���mm���Ԭ��0:ͅ�H�q~��������4��$���0hj����:`�G�8F�UŢ�2����L�wJO`E�>#f��l�S�=3�\v�]q��bn
(Y3�h���0x��q(0�:�]�YsO,�;�Q x��':�̦4�+�"x����2��g����������0�kW�j*�U-}TC,�J�'�a�?��ߎm�Z�x��`�i��أ:�Q`���:�\��4�o��cL���̷G �h�Ƣ�ԉ��t�Q^*�_���8'��O�텓iq�[�Pv�w*;����	M��O^ʿcI�<�)�[�  f���=�HW� N����F�! �kn���RE�/��*`��s�h�w&;�"=s%#L�� ('���Ԛ.�9��5��~����r����zmA)���؈��t�+��s�H����(e+XֈDg��#�#¢�@
�����"l/�y�D�� 	��KD���iG����ZG�~<T�/'�&nC����r������o+N<΂)���v!�7��9�� ,F�,��~9��߭Q#�]e��]ƈ��+-(4���.�B�d�[�V�K����_U�����m�w��b�z���h�<J�"��G�*U��`��p:��
䎋�jM���W�1S�J;\�����K�/�H������f�����}}�@�f]ʲ}(Y�;18�C����H䙞nf5��d&�5�aQ���9DUv�L���LA�W>w|�`�g�{H�HL��έ 
)d�M��gH���t~��]gRʖ�me��_�,b�����$^n���/�O^D�|0/��x�^�v(�!�Ti_���V�@�=���Љ�w��7�&iGI�ճ�W]��݁j1�����w���C���l�-��sбDU��P����,�=d��q݇[��;��jk;�������y?^!Ӷ�Yg����n/��$5--���)BrzK���f���;��{wML�k�z�{c�L\?��B�ǥ�
?�)�T�gG�S�{:\ %`��2��\_s)c`*Y��W� j��� !P.{���Ҕti	�<��Ҥ�1:����}���ј*>�LH;5�;�M��'ҹ����� a��I��O���{��Uw�}�-C:QO*-�댦��^Hm�=�=��!Z(��i�P��n7%�B0Ġ]_%v6z�Ǆݖ-e1��@0�zS�P�k ;�GH,ױےʾ�J����K�y�LF�fH.|.cMy�F�N0���m�&���S��F��*+~T|��H`��¬6%������Փ��� �a�g�@�O&���k�������d�e_uJr�W`�q�{{j� �v���ְ6['���{��m]��4�ԡ(� ��n�N^���|�1Ќ�I�o�o7֤32�i���UT�dٔd��A�L��� ���~`�	��	�Y1�?�s>T�����	pjD����,^k,t3ԧ�0�|W�\zY$6�m�%^O�6����AMwZ[�|7Bc{]����*
u'ɌZ� �0pswl����[�D���+�ԛ���+I�fj����>��g����_*�/?�Y��\]U�w6<f����-#�g1f�F���/��,���@�8a~�!G�HF�����J�e�S?1o��չd�u ���z��)�c�T��Aۢ�e��t�N|F���P�F컚�PQ�s�n��e��e�m�w����b;�L��N�Sસ5>��^=q�	.}��� ��-�5�����F�E7���f�'��^??N��8��)��::�;13w�ڰ��0(.Ä&�ۺPu�z1m
vu�!Dl/7�F8�6@�8�x�!�7_��tȀ��<,�e�+m�=xDX�M\�:�&Spط�m
|�y7�.�P�3�S ��DJY]��Ȋ �,,��#<����O�3��UƏtע��~�-K	���T��7?����t�o���#�s�y1���sYF0ct�u��
��O�Z�-h��>�y&�B�`:#SnY���ͯ����G�$���bq �PwF��(�z1�3FՋHY����C��f��,<��'��j�m���x���H�?ħ�7��N��_Ck!������~�E����c� N�1M��@���~�PD.�[��eњ��uC1KAi������ZW�߂�z�����H�oQ߄Y��2v��`��J��f)"�mLn0����J��if�`<���i|2Z�6�H6z�,J!?�Aؔ&zBW��(��pL���E�n�bY�o�p��iU�F��W�HD�T_h�KR�[�ԋ��,l����x��"G�_а��l�2fE\SX���^tC1�k{�-�X�Ŧ#[^�.4&v��ʴʓ��g}���5���pV� �Bw�"S�u���L� �0�W�]d�Iُ����Y�_���B�_���A���`�^����\R�����;��̲��Fp�+��h]�0�^=bQ�3	q�L�O��Q�R�����ڄ�y���خ+W�
: ��c���m6������ �}���\� #��/DP/f�q=���:Y嶴pa��7$�	�+\�ݘhm{�� �=�j��c�$��/��ξh����d2=�Z�th���)�lE!#��ڤTJ�vl��K�r�⇪ѹ����<��7,i�A9MO�k��Su�=����{'~�xOM� �w+��ޒ��W��wnU!��*)z��-��,�����P�$A��:�'�d^j�Tt�6}/k[Q^�9U;�|rY�&B�o΋i���҃Ex�]\�x�Y�ύlĺL+׭f����hg��t��(�՞陛(�79�G���:GEz=�m�h?��^z1�����I��:]��7i�-#�C���k��$X�B�~%��`K.U{��	��s�ãJ��L�n�I�M)ò,��r&��U��z-������j�܄����̓���OQ��&1i�����(��
�5��e�`c��+���¦�ZE�7��X�!�C Az����a��P���� G)�]�*o����绢��"�{�rkB|�N�C�lJ"���E��3|�WO�m�Ξ[�x�]+��*L���AS�}��W|9K
��=uB���W��նi�[����[�LFb�*�d�f����L@�R���g��o|Q~�����/�$2I�;l���[}fc���j�@�񬓍Z����	��B���|�wo��_,:S	���:~�8N�t�ֆ%hϘ���P��Ɓ��"Fg$�͎��~�H��kUL��e�!�l�����4��	��oq�U]��3+Ȣ��R�H�X8�Q|�����������ˈq�D��w�@Y�H0�~9��%�x��u>v��Ⴍ����+#�le�7I�w�b"�c��}+���KG2�fA}��}#��䶤�9J���މ�g�Q�qS�O���|�z�6+=g�e�͌ULϙ'E�GT,�C���ؕXK����гT1�M�!�5�_qp��}Yy���Rv	󧲓"�f-�1�Xؔ�{
�I�[7�_�|/u�ܱw/Z;�HjMhF0�T�_�^�':[&�v�D����}������Xg���Q^��H��u��	>��Ƀ����UޢG�n��dy]v�i�J#�%��k���a�K*iA9eS�]�5.�9 �`��m��0�7jKKI���ӷ��D�um�pX��m�Q.ܢIR"#���9ޱ�}w��^����3�����-|o���>��^��ǟ5�X���ce# $��=κ�NOoqiM�ŽYd���_7ӗȱ2A��xMC�ƴ8���Vv)V�X�)���n��6�J���:��:�1tl7��x޵����dZ��H�$X�UЏTb��$b���mU��T/b4�0������A��)D��
	h�GU4?�^5jI��e�f�L86lr�2�3یm�A��O�yk��,U��B�6�j�Z'}�5�Iq��)�FTL�>�3�rm�A)��9ϕЪ�tj�(F�:+��i-��n,��@0�6R�>�P�e����$zo�gJX��"%r`U��7o���z�g�YY=�ޠm����'d�NQ�j�aS�8���溃ɧNE!�!8$?�IeѶV�m{��eQ�E�EB 2�7Ĭ�D��a���Ih�Ĥ�^���Ǔ!�ӳ ��l���c�%D9͙�?�_��@㴭	眮6�a���Q�e�O����;�gL�C&���J�υ���z"� {AW�^�6�`#{t��,��J�[A�v��Oj��G-G^���<����v����vfi����t���fW�����4/�d����XY���@��6?"14v��e
�(��E��b�yxb�3��(j�%6����	(£�J���%ʯ)n�,�Y����wt�z���]x�2����'m�'���`�G=�$���u�zAn�A8;}��� =dLU@3�ÝĶl�AS@�8z�OT{I�s����j�����!��l�A��=Ñ��hw�T>�s_��9�o�9w8��f���to��۟�ޮ�
ѕ�D�}tJp;q�3���]���������F~%Gj�~�����p;�&ݻ�����'=����1�s�3	�>�n���]��L�	
yň*�5�rXO�^�����Ì}:�0�Ѿ`�ǆ���<�?��cX��_�S���`Wv�%�t�,bT�(~w[&]�F3p}�y��7���.��Fߐ�5Y���5��W�f
����./���KUCb����*`�/����%N�zycP(	"%`u"B7?9����U��U��H����@��c݉����9�_I��5�����P�3�x�g���]Ą�}�=%٥��fI�?����p�d��a�g���RRb��6a���AI�5D�<�����}�c�)J�su��z��\��U���12���4�4�5Z�o��=�ȥ��Q\��_.!��ٚ�83�uf���/ZX�e%��!3�����4�
�QKJ���b�����C0=:��i\L�<(\��rW˿<���o}��K�.<��ХRk����^%g�<�"�Gb/4 -��L�1���Gl����l���|I��tCBhs�D����:�ޝR�nD.��-1L�"]�2jbs�ӸUWC�����	"Nuk`�!Z"`����a~�{��6VX�ٺC�f�߂�nĪy���:s�׀�䛭q������~�*�4	�����Y�y6����5��ɂ����N���7	�V~��!}�/� �T�H����M�t�Bc��&�T�xCoo��w_2��K�fӠ�bK�J�\�*k��U��������x�M^lE�fyU�L �Ȳ�p���5��,TF�V�ȝ�At�ȑ�_t���8ƧD��:7�'�l��^ER{���61ݴ��
xɂ[���O\^���a��s�8ِ|j�s��4IF������nM����!�J��/��B��ض�L"��`���x%�6�R�r��8�>��J��X4��|�6��Kշ�y>��>�`)m�H=�o�ٮDD3E&���a�AQ�Z��RM����We�T-� �Dm٨�
Zi��٪�I6�򙒚K>>�3C��,�z�\q�rG���E�й}l�*u�Xo�xM/Os"2��� �,1�0���=-�՟� ���y"��r��)2���c	~$�eER��G�l]s̺���4�}��_YP����QonW�[y�"u�oԪ�jI��(8�*��"v$��G�G�t�M�]�}�-�l5�"��׆�D���Rq������.�������t�c_<��s���+����;4�|��3�ŽO��I��g^A�j�,0&mv LZ�2ݴ)����}���o����Ɋ���6�k��BXj&�������+)W��$�Kd����'$Z5����:�$���۲�mo���ͅ���l�7�aj|R�eu�ҹF���`�̀pj�mι8"��Q�Y�5+���t�i�r� i���&����O�G��gt�����-�ab���;ʣ۫F�A�Gmr	.�Ͷ�/�["5H=�'6�sO�%�Go�a�
�i������F�JbIG�ҵU��������@I��3�͊�ظy�E6 ��n|D�+]�+џЙ:�z2C�
��б���, �[4�M������ l������"��&vl����RH�P,a`Ot �ؼG�k�E~"�	�m�!���c�]0>�=�Er�y�w��P_݁F���j953�H09�	��Gin��du"Jఔ�7����]A�o=��-��>B3�H����a�@ �V�Da��l�iq�}�K+��P�i#&�Χ4S���Bw�H�;�m�1��2��gu�]�o���cr�$��=\�f��l
�ϡ2�!�
��w�S&�/�<�}��?�9��s��^���6��n�7�+m!Sy��������{�!�AI�4�4�I�QL���R3� 6�kϓ�^P��D��Ps��;�N��7Gf�s/	>�&�9EFVon3Uj�4��sE�@;��O����s���n��r�W� )}���8e�R/@~�Pr�\;�`�_<
�D��踨��I�q����X�).T�I�1`�Q�%
yL�#ڞ�XG)oy`/_�=�k�=\R+&�l'R����U�[���kp\К{�oo`�{S�}%C�)��w�M��D����3G�������qW�ӹ�$�"vì92�?�󯞰��t�O^6k��17�v'|pO��æ����������b���4���8�u!�3P?R�l�;*|��*�<iN娝��{>F��{NI�0��t�2hY�_?T~�W���λ1	����ha������jJ��C��`u��� ���j�.t\�W��OBP�|J��N�����k������Y����Ac��f穿�b�3����z��GS#�±~�B�1ݷ��s�U`@-y�{�o%�2A���0�[��_��t���7`͘���#�]0t�����Cl�wS����4䫶$�<��j�0����ؿ��ǼQ��:Nώ���d[�';}c�b�q ��h/�rz�"��DOѸĜ�JԽ�}�'#\$��%��H��MYL��+�;�	����L���D�������v3���3W��({�i[$�8�v?h|� -�*, ���"�
��-6��Y�iEL�ͽ���,�<��ʏ�O��Ϛ[���KI�$�ٱ�Rh��E�=����Nv������2�G�B&F�!���� �y��wr�Z��֒1�������OE0���*:�v(
��,!��VX�19��=�%�}�8���e�5�,l>�pqv��\e�2]kn�����y���3�t��&�C�!�Y�1\��Xy�%��t�0��fm��uᘧ�:B���DHUí���l�z�T�%2
�qqXTK�芅�CzN�	��a;6<Yp7%�s���wv��s��#FP�P~5a.�Hb�e�i���.;hE�E�*BucѤ�2f�L�/`��,*��+����X���	�%Lf��3��ؼ�MgG;�^q���R����)���.�@�<*��Χx��ŉ		,�Ś��bgSg�0A��563���b�?7�h4c�TI[l"<�ku��=�X�b�۵�M����r(V�6r/���c��V���'��.zl=2��u�.���@1F�gtd�O;�.�qI���!,���a0aF�ujcd�(8�[ɢA��!��Y�$���P�$w��Xa_�%��WU������i��_�ˁ-��E5�i4�8��b��z��q��.A�m�.ő�p�J^�¤�y&��sb��kbv$��=�9�C��(��QaԔ�|��6�)�1��j�2���7$�2x�bkO^���e�@.7lGTٕ�f#藙�0�sS�I�e-/ھ�|T���$��!�c�h���2_U��"ʙ`���n.`P��ὍD������Ij/)ɵ\W,��\��D�t��q���j6�*F�V����{~��p�fLz�v�p�����&�,wJ<��b������_�s�+5��H�8���b�G�,�~�LD���;����8>�K����#�
���Ew
�߅�����s�`,_�Q	qɅ'�>ǐ�]�P�f(D���q�A(������9�-�d�wn��`�7��`3X��Sn��`�����4p-�#��rmYWO���!���E��B�gp�-&�����a2˿Ca,b"�@k"��]搼�O:��O}D�0���6a��$B+b�V�>y"�����>���j�Y|�,1nZ������~W��Ꝇ�9�B=m�~���� ��F�	��3e����V�Ey#`�HZ2�!|�]M�E����]�֋ �����mqn�Zx��������h��[gj~d�!���Q�2��[��}k�f���Tݽ+�Yp������o6.��K&
�;f�~�VH��-���B�cc��E3�8N�����I3����a�[�@R�?���J��3���{hO�.+�aӐ�0�Sݲ̍�Q�;J�x���ىS���4>V
��r����8;s)CB���V�́;Q�]��=���w=��i]��c#�[�E��<�߹S�Ǘ|}��eX�Y'��Vk���2rYh~b�vl��m�Ԙ�*Q��l��8ʜ� 4-c�oW���`{]�F)�����Wv=7�?��d%�\4�J�&�W[���XZ���oiRQ�+Mw����[F�/P�P�L%I)��0}�,䖲�v��.X'���k���:+h`}T~��/�0car@>#@B`ie�y��5.�� 6��h3����٠&S7�s5܉W���W�d�Ie�V�� ��o��c�`(Y�^��l����K����a}y�J{�$�4^���o�W1aLjw�&ϛ��a|���"k�V� �@��������8t��݉S+�ꐁ�C'@���s�ݒR��o'�,oWdP�
���[�,��|!�[d^��q򎮴0���h}V���)[O.��>? ��������*i	���K>K�|e:z��!W.�Ք���~[lN;ݬH׋�]�c5�s���*�N;clJP������[�u�2���]ԙ��O�@?���;f�Go�B�F��q��Ck3���1~�o_��
�)"w��L��J����"I�n���[��à6���:�Ow�c*PT���h|�I��|�*��ld��b�ި'��S%1�L�����9�'��l+�P�}Te��϶�A���SU����|ڊ�I�I~}��s���3�U@�����_��d6N/)�`��&�@d�]�&��]�F��S��=@�%F�F�ٜ]F�yI�����ƍ�US��V�U�_������*l����s��b�K�4PX��=~JX �5_����'�1V7_�c+�F�u.:�����}F�g@�{ﰂ���k��f"�Bh{{@)��������T�5��Т��j�O�ʬr[$
�K>�a\�L��޵߷��s�f�$��D���uk���(�N۔e8a�x�F_+����iڱ}e�=t���*Q��A��#W��I
�w�/-�
6q�D�|��H8�r���U�6�q���<��=�ϒT��@T�ES|j]��n7]jo�;���ń���ń1Մ�TECx:�sOęV�+#��0��Tn����+m,K�JA0��7�փ:xU~�nK� �E�= s3�$IW������G�z�������Ƴu/�Ӣ��e���X�6��O��(a�z^Te���a��?�-��N�˭W�ht*߈�"w��\��� �
r���KBe���چ��Y��>%\k�y�O�hu._�td*�~a�����Q�	�Ak:�s�ks;R���p(�^SCٱ^� zp��v�↷]�����ũ)��L�'����gh�֚t��Q]��G��.bV#�]�K{V�u�>N+G\37��Wa��̚�GG�n�Wo�_��1�]=a�w�����"`]�k���G��B��.=�N@�6^˻A�ǒ�k��Ti����mP�R�e����'d9x�f�v��c9�����F�VxLΓ���{����E{_�Ma�Jﱩt ��4q	�@[�,X�0g�z�H�`Y���w8&���Og1����5rK�$�rӓ�f�,xB�|s��{����tL)�7���K��<�T��|��iM� ON6������T�x8,��袉,P�6*t��J��-��"]'�x${�h9�H��#u[��͍��)N۸үr���ϙ��ۘi�1a��]��e��W��I,��-��Qݒy7����/���f͒�r�%�U�?�Q��� �S�3)4*��#���Ø��u�L(�[����S��|��^.;zd�]y�/�Sɉ�kSO�����Q�߿@Q�c���&xz��l�ey*�j��syRb��Eɳ��˲}�ƋZ����8���n'9]��͡������`4B%A#(�I�J|�	��.��T�Y̳�k��0�.��Տ;X�ѥ�ȍ@��O�ض����
�
��\Mq�X�w"�F]S��m�jU�8@AuϞ,Q%�����9��Kט ���Tv��u��0�EҴ �S�Gb{�(��ZY;��{�\1ؒ�L�s(}s7`�dY�o��t�;���Wƽ��s�6�q���f��������Y�r��7�H�.��n���b�+P�M���ݘ�Z���E�u�*�s�d�jTWD*�W���[�fΜ'�f�'���F�:5����a7,�^���D���D�!��{8����!�H@���a�lN/{Ζ�������A̗S'��rf�mlg��:�%je� ��X�9+��du�#���o�k�a
l�R��U��B'o�x�j�-d �L�^ ���8�>���.�#v�X�1^�b�P	۽WZ�tu^����8��23�!�B��rrMc�8�������B��W5���4c�yFeb7
=b���!u�06��t4�)�J������,=�)�x}U�Ȧ�S��JI�o��F�B�,sݼ]���l� �K�t�H�Ǣ�������t���|ҬK��T8 �bBOq�0��*G#�s?��+���7j�)�i391�ar��r��Z���')��5����������7X��w�hd|ڍA,݌Q
hV�A����S�A��C�Q6�5�1�~�H%��"���s�״Gh��EN3͓�G�[��'�4a�Y$-��X�X�����B�.���;|c����*���[�
]Vjm�m��a�ϕ����"��\���_L��O���9����X���,#�f�Q>3Ybg�
>Q��@������A�	o@�y�ܸ�Ʀ�TW6W�"�q򸒻��4H�F��d���Nk��C�O�����S��,IH)�[fU`�z�����[�Q2[�1/j~:N�C�r�8��1�ר��TKc�jl�ß��g�as��LxK�\���$��,<Vg`��*�S=�U�(�m?Ì���E;��H�m�O�H� "���Qf�w��Bs���H������ޖ�|�u�0.7���9qT�C�z�ē+�q�*U?�Cw�����:Jq�;���s}$ʂf]UB�E�#J�n��NI�Y�q�������՘ ��>p��i�)]��C�G�76/�K W�v
�h��cX�`�E�P`��
��˄�D�>(6rZMS�9�|��8F()�J�YE6���E���%�3� �qS�i5	*�m�K�{��v��}�f����'��%����;%Z�
���?�y�}6B2t-���9�Ά&Vt���am�v`_���..�VVh�E*�J� <�UG	
��Fa [�����ϋ����qg-nb+ėo��Wt����Џ�Z�Awԑi{�4WDp�r ֥�C0a�?6�lY�\�[�S���$�{z�-ݓ�CDo�cRy� �	���~J#��&��z-��ԑK��8/V�#x�M��RxU�ܖK�Z��{�eUԄ��V�0,�3�_	t��(Z�bȍ��K���4��́iQ�ك�쳿�o�������>�Q�K�D�#����a�"��z��e[�)���j�n����\:�ᤐV���8�~72�(��[����(��	�M�n��$+���p�
`u��h�Gq�r�a{Yꂼ��z�շ��1X�

�����%�]��dU�)�;fG<� S��L���@�nU����u�my�~&D�}�Ң�
?E� �I��9����^�muNѤnw��4�q�u�
V��g�	���k�h)fRGzZ@V�����NC(��� E��F���Κ���{4|p���mNr�w���E�Q��b)/�V{�+�ț%��S�z[��nrڡ j�-�����"���[���NE�E��ߕ=q9f��M ooIxM��l9o�����iQ��Q���sg4�#N
�v��縌�䄒���������܏B���h�
K�M����gZx��đh��eT��:F��ؚ*����Z;�/�_c9$wH�ÓY��p�W�W7X�2�a+���S��ڦFA���B0������ o�ʻ�5JgJ����Uϭ���H�v�R6�eP��߀�<�i(뎶:/pΛh3 �Ϩ����<��&�)���P�q�$d�M_�[R۳vs�n���G-��F�����_Khzݦ��F��&7W����wV*k��u���t���rP{}���j�����Qn?Z�?�R�4�e�&΀���b1y��39�Jr�U-���+xb�j�<�^���x��ړ�G���hY5]?j֣$�!���s��N�W+�Ƥt���E��GU��}
m��
�h�B�`���b$r�&�{.Ċ�{�$��1�,�!奂
�ɓ�TY<z][�U��~���Aï��3��\��<���J���H��7�D�Q���xbE��F)H� ɖ��J�J�����_�sl�z�U~vS���xCH��e>P`<��w3)�s4#��.Idq��H7�R�3��.Kz�<�(ioV+����$�S_6���nQ����_�ݤ�S4.���Ż7?��_n���i���,n���tUX�d :��lFm����R�s��ѵ!����4(i�Y �k�ڕ�Z�d5���V�~yx�X=�o�7)g�Q�r�����u�$$��z�� �A�#i+\�w�	Y��?�0�#/M4��:����r�s���U�[�@4|��ɪ��w����zFI���5&�j ��A ��Gֳ�&�6xz��vB�k�KK���\�7
-���1���\0G7�Ś��cL0��3���F]���̏������`.6Ɨۗ���O��K><b�>��w��d�;��y�[D��.�#�)&�x����Y�2������(����s5�D���Ⱦ���b�y�̂%�Ziu��tr���e�/[���+�X撋-O��'o��]�M&V�1]���;�.nm?D!u����������RU� &������?�E������bҨخ��Tk��(����劄4%5��W���B�È)�8��В�����Ԍ+�?�b_��r/&MK8���a�^6~`W	�z؊������K��ָ���?��u��=�z(�o/��L�LV l͖'o�y��|qг���M K���\�!M@Ʋ{��ԑ٭ˍ�D���X��v�2�t��}\wN��[�l6�8����� �����ҳ3�7�#D^�J'd˓haS����2�{��k���'�9g%|D�[� �5e�h�1��k�rf\�CI�����z�T=���q��-�gѨ=g�0���Bj�G��n�T�e��R+;Iꂼ����!}��coԇs⾷ߌ��n/���׋j9wt@��dv+�[1��
�o�𶤋F�s6i	�*�[�AKk ne�>�F��,vS��{�i���T`h'@��m�GBע�l~i�����M���+)��PC¬��(��8k�9m:��ޟz�>	�ç%�r�~*.H���yp����1J>�e��mp��������SE��$��)iP$���O.V~7F�+1i/��d)�m�5�Q�V��W�z��\ˢ�����|���L�btR�5�z���x<������lDI�g��;]���I�8�f�U�~��|�9�<����N3�s,9�^@�P���J�Ro�MI	�r��!OA���Wm+������NI+ż���<bs���H�B�����ȿ�.�b�7_Ec�Q�8������H��+>[Pn<x����m\_ٽF���<���,��i�/����/�Q�
Jw�;�P��{�U��>�t��+p|C�M/Oe+����ؘ����~��>G@�����e�^ʌ�Աb�]��������5y�\��B"E��,�[�jC�0��`���O�C�������Ƃ�ѯ�d�C`�#;3�PVSR��'[����_��\���E��om�t�̄\�\M\Pa��K��Xn���⇥���.u �X|"�ܶy���Y��N����4�Q�Jx9�:�
c�e]f�e�]��"ZT$7�_���ہ_�Dr����3mO5����2�{=f3�k�-�+pM��ũ�0����[z!o���0@ԁ��a�ߓ��i�3��������u�w�F��?�D.H�@�w�҃��2>������F5��a����~n>��WE$�i��������?��KίS[6H�(��v��Gf���8�� �hk�\�#�3 ~p�eR�X�� ������x42��;U����3ֆt"s���=�h��E$�)q~��2�S.>Ǎ�����3��2p�b(P'�b��d�lqϩ��|9]݈�q}��Īc�mQ�ք|�Kg��j"-�$��o/�&�H��"���kɑ���:\�ᤔMr|��+T8yU~�]ѮR_�z�C�_QX�5e�)���=�aC�TT�B��YR��85��)���fk�d�:V��W�r��^`,Z�X�G��؋���V%�.9���h���vj'�f ���)�sф)k�{9vB��vR��T����� ��_�������2h9Ű?^|��S%O��f���3��u"{��e�C�E'�}��&ɥ/[����KU��Y��"K�"�x ,e(�-.)7�#��M�*�� ��w��`���������=�e��,�'S�.i���h�7�g�=ӗ�NM҃�0�DC���yئj|r�%�H+X�)�dZ@3N�-֙�C�P�<Uc)�k8V7&�P2�ym�^�W���;�.�?r��� R)�o�����]Ƀ8��� :�Z�.;�]=�-���wA�_��ETGKWS��AH|�� ��"o�*kk�mV`uQ���AQ'4�B��ah��~������l�����h��U���i� qZ�u-̃7�c�f�$q!��H�=�ClH�|M��
j�"����ę@�s���y�V��|��/P��:̨��I_?��*1��RШ���eB8 �iQ��<C�X[6�^���G����F#Eƫ^�2<���,7f�@?rӦ����.:�0v��Jz%��� lh��)���Ǡ�K ��j��"�k����$���g4���0}��_���s�=��,�x�t���������=�u�������à��E�����<0DJ���gL8����?=T2�!b��SC3�г����Fi@�SGKٓjH�Xi�p�2�~=1½{�\����:��{l�#�o�½�n��9����%p��"�]SS	<G�����v%�f�m�mܨtp��v�M�.�À�X�	��F̔�q�6k���D
����CBʩ��5ܐ)5�.�Vmb
�:���<!���b��o�_���r*�t�i�!ї�7S�}y��� ����4���l<�r�9߅g��!|MW�� >��sI^�o:�܈;䧥8��d��`�,�ccz��-�� �8v��+��j2g�ŖR���ْ�����nz���o���թL�{�1L���hw<��y&�� ��f���޼FQ�+	�kl�v h���+/�/�lѹd������3'E��p쫁�K���f�s�<�㔶��g�BGI�?�����]��8_�6`��ʲ%\q�8�Pg	��;� k��K��>V���r32E����y��%)�ԩ�6�QkF����.0}�w�"��Ns۲.�w�1F6+�
��EIk::9Z!?��5�-3$²���R�u�6@�ءk��E�w�6
��(���M6f�J��"��~bq!�EV��.��%����<q�ݰ%mq�/V��so��&� &�1�-N�߿����2����Q};��ګ��I���՝h7�W �T�_FZg���;�Kƿ�D5�_#�o��#a��I��2�#TV�ɳ��:q`_�����Q�Q�g����i��bjU��WW��P-}&C�^�/�F;�K�P�K��"���}�R�Vm�ge
#��p�����!��t��⡎S�x�y�7Yo#��ahk�5Շ{r����m�Y2c2сq�a�����BȌ���m���~о�c~t����r����F.�{9��:�_M��@�EU~���T�.�;M�!)*�ǌf>�,>2��K�b��)��hq��*�)Y0�n�!.b�����߷��oz�+���7�AN�OUH�uϴ�f���a�,�jM�B\�9�%�R��N�L�DzZ�,[Y��m�<�ą�!*#���ٳ�â�K��d�����m���>��G S���q�:�@"����˞j�ҏ���+��*�g}T0���r��a��f$�%�\��SUR��A�,�|���8���F�4zT�Nc3YtNǦq>�ߵ�=5k��U���ZU;n$����4�Nh���C!u�}t���<�1av�u8Lf���1���Ɯ4� )
���:��k[���D'L}G�j��z�~V'l��'QE�*wpi_�m�� ��9;�a�q�5lzSe���"��Z���S(�[癴c&Kp�;�����>���*j�٤�;�����f������R�pt�JC�re�9DǠ��[��,�*zټy<3��
�m.a����]����/XAa1�o5̦��eQrq���l�a�bS Ƶ��P�8r�z��&�I�+"�V4W?5[\��W�����m�e/����n�ͻ��e|l��9�;����QA�����3�����~�jR)AT��yp�L�E?R�a�(3�~���?�3.��@�"�R����[�u���n�����(���K�h�&���
���z|�����K3xZEUS)Z���VB;�e�y&(p�c]e͝C;��0G���Es��_Z!����RO�˸}��Wf.� �!f�_�xO_��/�3�rNj�D��e�{N��b ���'�^c(�+#�I�[T��������w�CkO��5�%YUn����hJ��l�y��Z�j"��9/��b(�8��p5��_�$\9Ɩ�%�W)&���X��fo�A��tc�)���R�	:�������+��U�Y�GEr�Ov��W��i�J�����r��@�Tk��d��J��f��c�:��a�Z�X�$�����yu�&��&��Bs����I"��'�.�o������=�.����khޮ�Zg)z�܍��z��g�k�-��x%�2���TAd�$��G���.���1m�!���I1W���<D�C�*}��6�I4�^7�@��F	:2٭ܿ��7�S:8�����6詚2gI���rS�ݥ��J+�Z��ZF=���tx	�1�l`T,��toM�	��^p��Dv��K�d���LKY:�*1�/�н���,B�;��[�ӝ�֭��ͦ���}��1�<�"��2Qz�.�����f|�i�!q�/ :k���r��oWc��.���x�õ6��P���t��bi=zL�ꛠ�<?�r |��Ȫz�A��_��@rc<���v+�{Yψ�.0ۅ<alv�Q�)y%�[�w^.�'�K��� ��+ѧ?�G�:���m�p�5���^��3=��M;���~3��#�A�*]_o)���;BR�>^XH��y�/��dW��A�m��/���4#/���
�q��)�g�A�YB�]�wN�5��m�Xi�ţ<C�m��6�ޏL��K�e�]�Xz�bZ��U�ΌͰ�k^"��N� ��jj;޹�=f�|e9�҉Ml�T�a�W813���o&Ά[��ZJ� ��8�?�F�[���� �DRYʇ��������@��9�i�z9�	���]k��6��Mu�w�����Ũ;)"4�E�O&��>K�S����*r,�
M<0VN �M�q��DFi��M��	��w�
��U7� X1��ʆN9"�� �����	i�WT�W_#��P�� �8�p{	����1.+-x���a'�z�o=�����p��8��&��]�Q	������|-�a:��nH�	�������뷚6��nm�R�8�#�$@�azC���7�'(7=��n�a(��.n�
_��O|%ç^�T��ѻ���f)v�o�pkA�GBF�\��j�x���B.P*kz!�6������U�O3���L�pR@��WD�I��@��{�D��	pB"%���4����z�?��NgB��ÜB��\q��B��63��?���j�)��)�WU\���bH�����B>�������!�O~������>�E���ճ�(���>�7#Xq��+4��Ӡ+�,N�[J�sh[e?�-�bӈz�������u�N�Ԓ>�[�V���Sf^�u�졇�d�{�ꊩ��P�W95L��I�
{����V��� �Uq��Ӆ����e���E�a��WY�j.��"����C���>��:�.%�x"MS���,4��g��pD�%#]"���^v>�{���(�4�͂t}=������v+��"�W;8�|<���ý"����.�v�=Ez���0RQ.^�t����f7pO���Asg���o���x,ϤG�6��?i:FV�ݥ3�{B��cl�џ엜���VL%�G��t��W�J��<���F�RC�3�${lU�he��0�m���|%�nhZq��e?��^U!u�]Q������߀�R_5�3�N�+�:���� b����7���U���EC�èq"{
2H�p'j'���ݪ�f�(T��{$���`@�"�,C��a�1'�����*��i���w:���YaD�5v&vn]N�_�,��e���5��:XFm�M_]��l���r�;�,����{Bɇ1��n�i��gT����(:`�o�.g =�3P������Ξ.g����(bR������|?���$5O�Tma����d9��F�+N�����>���uv	N��D�s�V���y�\�E��U�H�V�U�W�1���D��
�AU�nX��9Ǯ���/F�+2�o��J�J���ww�՗k�<�haRcE`X�KwL�͊ＤG��r�m7#ʚT�����zq����L���TN����q�S��A��l���;N=X��j��C��\�L�|U�o����lv��)�kB�::��j�ߧ�M�m/�d^��������1ʚl�g�2U�Zys��-��1�9C�0@S��r��X�	�Ԅꯄ��7�����|p�g��-{���qz{�1KÊ����n�����p�J!�g����w�f�[>���+<�z���Lp�=�|PZ;,��b��s�H�����ݺ����V�7y��rK���Tw��2�x1E�,�\ĩ���$�!k����/n�Ѽ�R��~�z�Q{<þ����H��m��H���m|[UZ��sι7�ZT���V>R�|G�����g��B��Z,q8��RR�Ŭ-�ds�fS���/�U�Z����t�l�y���v��2K���N϶Kh ���`�YZ��5c�����!�@�T:^������^�BFtl\���ya
�`�_N��V}�[��{���Q@�w�o�j5�O�O#��	g�79�!�-��Òk�W���p�px�
<���|,�\�)�X�BU�=c>���$2vn1���Ǣ͡ƅ���#Y�ο�i���`f��;gF�5��w�i�;\�x��Cnw�Ȣst�Ī:�$�4�����\6P^�H�@�-]�=\�pJ�(}/((4�{�vo����*ii)�9)|-�wP��۾��o4ԙ�t�.���C�����P�B#R!���֒��UU�v@t�_��7m�6��-v�@S@3�)�神�pi %C��|�T9^P��k�%�����cI��[W�(m飈��03]!��J��!_b(X�j�O]˷;�%�t�c&�S�%dgu�yѼ��r����op���$�A7�v5�Pm���2�#x�WQGa�l��������uS@��4��f��~�<ijoE�՝l�]���A�����t�̽B�M�̡��aEH`��ra+�u��/���'���@�mp&�O�L�Ype��D��ɣx�QsZ��8��3�HR�� ��ُ�&�@�JP�.�TT!�!��+F3�b����x�B9�G�_�?�+�w���@������$	�B���f�
h�Zr��2�}����G��X)��يmSQv��-e��N�����Σ�?V]W;��&H�xC���`�q�W&6[�w�(���r)�+YuZ���^O��R:x�E�)�]\?�/��kj��z�1�h�=���8���B�
��`����=C2H�U� =9�J9_[t[��%���低!���٣�/(Bw�R�߶Z��Ϛ��z_�&��/+�] �Pu�k�܇���%<�ռ��Nt��dO˲P����f�6э�!�OX�΂�r��y���"���}C㷈-pe��0'~e�q)���1ѧ�ޚG�v�X��&�n��"xL�i�i��XW�~9e"@�؝ǽ]��u�T¾�k�u�7��=�d�@<��C�<�s�z�6���-o-��Qzu���h�u��ykP�T0� _�v5�Ζ�����\�W����j�نYw�Z������D�{jrn�׏��+=va�� :�U�a�x	6ɯMn���܈�q���/A��dг�屷�*�cX�@0(wM
4	�_�(��F|o�h
V�&��ɂ���f�����Z��g�n���\Vls��XH�#ɜ(�N��VJm�jm�r������9J_BGA5;C�!}��b�B|L�2Z�h7i*?���
�/H5�L
�����r;�	�~����+ל��5C@��A�9�|]C:]� }� Ц�xՊVd�4��ǰM>�"I�)z�hOC�`%IqcѨ���yA~lo�h�Z�=(;v��7��Km��!8=�)�𖟩1��AYR�QDc�V��o�����$N6N"7잸�@��1\ �#�R�KPڄ�d��Q�Y����
��xHw�	�U�G[�/�[ �̫DK�ð5oV�qQ�I�x��Va�	Z!d����'4��?"n춝��b�/�%2{������}��:)�_�]F{�nOǚb&j��{���X_��ep����U�3灂>!�tq��!�����Zt���Q�^�-t<��b	��ju�}��;��W���1ʓ󮏗��ghIf��<w�bDk���4�/�4`�iX������E&�pH�e*k\9����v�/i��9�g��*۔h�87]����@�!х�t�y�j�ۮ1�m�^2[͜��H���R��,��;�2�K*0R��1�	p�̺����3�#�2���i7��|
M���-���K���<j9�k6ò����'�ʾ0J�C? _=�p���ޚ��ɘ2�R^��@Lƒ>��ϼlɛ�Le�|7��'�'���D��&Y(.�>Cme�Ӆ.oPZ��3�	���c\���z�؊�˿F��� l�&׳�SgZs7�t��P	��-�VP����j��(Fu�J�V�G;I���mb�ύQk�n�-�B���^�IN �J�L�0�||F��$�a��x���xV;�1A�� ǳ_8(qt(�u����Ne4-�����d%�p��dl��b���.L�h]�\�k������*�8s�>�y�IQNd�m��v�{_��<}.t�b�k�	"�@�N�L#йK'�Nx����j��pBN�uX��`ݐ��Nxā� P�8UNސp>�?~�
J|rc�U��S���+aN$(���ꘃ���5�J��4�{��7Q/�G��N����D�����)(�˓s�Z�ڋ4�'�5�A|���L�V	���t�`�֗��M	S�E1�=s1�v�����f.�s��I��Ǹ�z8CϦ�|u�f���	�F̵H�+3��Mm�[_�9��3�N�
�������hM��sT���l�q��&�Gx�쯯&�`Z��1�_/+�x8�y[��B���͵+�����^�����)�~���_O���;x���7v,X���@��PBˊk�u��4Q1�۸~�lo�Y��[���t9�'s�vc�5�L���cg�g!��.���Z��yv,`�OvHEi�S-�����,�qlޤ�(����㓼U�Ш *���(��I�5Tma�T%�8�'�MI�m���a�O�m�Ž����׮�|�cr�m�f���j.?W���(�&Z,�/�� Ѩ�sޣ���6�tgd���9��_v�1��~D��4��e;�%�g��-d��DL�(�$�F�ajq��5���s�%sZU�P=���c�[���{��@)쎬�;Țo=��9�D�V��]�	��|�|�R��n�W�:ͻm�YF�Ȟ�-��#���t�[E�������؃������ER��b���$��V��۫��$P�|O\X������+Ѐ�r��� �ٰ��wL	������'�o������0=�t��n��gNI��Ru��ut.K���Ǭ��4b.) j�g��ώ�}��g�Z�r�|\�3d�g���M�t�z�wa�E���J�oT���=��w����r���t�T���L��m3B宲�L�r�*��Q;|]����&��2oT�e@�<���R �󵁵��%�YE0%^�Q���R2)H���L��Y���cm43�|H(�|�?�\�qͶ�����Y�>P�d���3���\��r��F�1��z32s)c�)�ԧ�)��]��8By�sl�����>Z�h^}�U���/O�粵p������#2�ȗ%�6M����Ξ�⅔,��ơ�����UG�7�7]"���&�0�h�)� ������6��9�p?e�3��,�����ѱUHA?���[_ɿR��|,b5t�CD��.R}�K^�E�{?������}���<�*x�bp��!E�4��G.ʥ"5Y���t.�O�l�N?�y]�w��}�ˇ �4��6|2O�
U*��7�>�������t�'��}ՈEE�6A{��V(6������t�D�`n�~��n�o!�}�'�'�Թ<�����o����� :Bt�}�u�!K��j!!���[9��G���1ީߗ}ǻ���ԥ$�I��O���2���|���o�>�Wߞ}Z�#E3�E��nMS�5Ӝ	����<�������BNȫ�Ȑ�.
������t�~z��]���_�H%��f� �Cm��#�.�Z�|E~�WTJ���䆈"l4I�,lS��n���u_����{�z�=g�lQ-�BL��L�_��P�x����q	�|sG.$�Zy�R'��k#x�=0Wu/��O.��;�e�}!�W(T�F�z�A�~��;��PШ"�<䴗�R��T]6Af�q�pn/���ܶd4ħ��3�u�p�=��z���	� /X¿G����!����9���?�n�vQN"�l� ��K�9��c�E���{@Ey�L��kYk�X!����H��q��i�U�k�6�b�J��,���̻T�]���t䥬�Dnz��_� �ٱH�.�?I�~~v�qx<��ОV���ހ�����C�
�:ܤ4w����T�j���_�OL6���g ¦�2�]���?�[�����ǖ�(�h,6U�k�b.l�Ax���4�R��J�܊lpV���wU+^�����u�ԗ���Pن�Sc��(�!���An5�]Z�Hw�g<����#�[2ް�n�UF\��O�5Exe�g#Np��+�F�8g�Gr۱?Pjy"����^ܠ�`�s$��\��o\~j	�k���9B���'���ͽ�� �l��u��.�����mv�=��yZs�7,:�]�=��j4;���� ��˾�>��D}ۼܥ�髏c�7����*ev`Y�?r`�L\ʪ�R��7Ų\H?�F�4�4�r% EA\����P4~�����Tē�wut	h��{��C���O�3��?s�2�&
;���BH;��:V���N	c�2�߰�aBx�+����O�o���) �%l�pT���Ȓ�>�=kmα���.�O���Rc��a���D���`4��*�Ed��I�r�^tN����|TY�+�$;��������?IRU<�[��s~zW-�)�X�[=:�Uh^����l����:�@ʦT�o������vT`Y�8@*��P�q_��
��I��y�F��IeG��P/o��b�q�ԥ���/%N|熷�F�;����2����B[�(�zM�zjg÷s��w�P���ݔw�0�.�t'��"`���������N�:�!��l�p��vM$�huw�U����}(Ӭr0oY��ux�M��gP�˲�D��Rʬ|��
����ukP<���*6��y!CZ�K����MP`�h P��&��紨D�b7��?�\�3y��w�m2J�>�� h�����8:
5wz�K���s"ۂ8qFSp~j(�j<��9uK3`��r=}F��\��w����wi�l�]JZv��PQ{!u}i�a+�'�W!H�
p��vW���{�4�d���rm�6@Wu���60a�.��[��a��_��)7����7zw��9���`[�@*��*��ܗC|���,P$ap����/&'#g�1�*��WƓʾ���|�k�h�L^�����E�� ����(zT���n�w|���>攑1�09�~ۖ��y&ޔ�A��]<r�*<���+�o*�r�E�ɡ���0��^1M	��飾��!��7��}`* *Q��2�9/��@Y�g$��-��(5Y��AN{���λ����{gy�YsSֻ����o���.`����9���BggFY��ˉ���&mc�.�\TJ�_��B��5��W�J����t52X�Πw����H��i_�7B7{e#jmhtTO�8܎{��l,-��������i�gٿ��l9�����o%x��|���<;��m�O��+"w,C[+	:����ѝ�SU��e��#���x|�Ms�b���Bk=3�Re	4ʝ}nE��:��s��/� BS�T }�U��CA��ĻN�Fu_6u�+)� ��m��%9R�&S����K>C��{G�� UD���ƱA�>�{���a��s{������h�,��DB5Ycrz�F����_�\+��:v�Y�����U],���E��\�D|�����ЁJ낺��Gr�J�f���޲��C"y~��e��F~v�P�8�~��]������*}�Q�~�ʡv�mңȮ�(tiL��s�K*���*�<'E��	S��2]q�~Gk�_4�ۗ�%�Ɩش�;����b"�6J��M���&��H>Z �hZnW��%>��J;���8��]�Ҹ�V�w�:Y��3�d��ȕ��joTH��I/�����2	���qs�b!���P�ʹ�t�e�CJ+�����Yiب=X��s�c�Aքah�^��[�$Y%�!��I7N%�{ySt�dG�{֐���_*�0ӿ�7��P��#OU	x����N$����K�1B���:��Q~�5�v|kh@hɭ��y�6r�o��۳#�����I} �}-�O_�&֗�N�l����)�ξ���%�6Ϸz��k���j���l��Y���X�5Cw���N�(�R�+�/ x�< ���e�ޕ��������dh�v�7��ª�53������-J�=&_���$
������>�oL8G�a���n>�3���L0�\)��@A�h�������\��j���m�#e���TA�R��1��`$`����\vESYsI�2(���H*ߘ���'
���EǢ�S����a��m6��f�/Y����XaBwZ�7C���G�d~,v��@�(Ɗ�ڭ@��K�Įm���b�HEu��&F�n���k�`����S�Q1pp&3-W�o�����C܎n�'�$�Se��_���lg䳙���,�5�H] F�a�����«���0�F}���X��,lB�i[�t���Q�Ȧm/ʖ�q~�rI���D%L��1k�UE(`�Ί���԰X��V\�Uv�$�;?�JwV�^R�C�g��R�p�����������MB{��0�_Ľf-�v��~0B�I���8�X�R��l�V�w�uG�^��}�uy!���a�lВ����f�t����P)&�ۡ�F_;]g�I�a�B82K��{�-m���)�E�;:C.�A�
2�]K^���͈(��V_ȘM�#�>�@�B_1�b���7X:(��t,*qĆ�I�֗��G��z��PH��*�����[ !�%�4o`*�O\�XI)�����:�شG.�T��pcM����+�]�0fa߾�Ƚ-�S�����6��(�b���Ӡ���
5��6����|��٣0{)�uK������_ʸ�rƩ��fݏ�(a��q���[���8����|wS�䂪Crm�F!K���y����γtFN�$�l�!�覇��;��G���Xֳ�&}���V$i���_tp���VU�����t�l���ę���D����˰�(��L$mѺ��-^���uu�_�RQn����G[%Q�誻�)<���� �gGXACq|�KJ~��Gm��C�]�� j���%uG���	�׺H*/>�0�� �$���_=R��/���z���L���:��=v�R��is^&�<��b|.�θ���wmC�;����@#uk�S�%���y��l�b!"�����\�8}�@HY&����h%��g��Q��+oE3���ʀ,��z��Bn�SUl_�`��ї�p�q�n}zN$�� v@��:�i��F�*�.[t�k%�,��3��G� +8=*�ᾢ�Fݘ�
�F��K�$ƣ����9��G3��SB�\��sh�;�?�9ܳZ�m��?D����6�'�t�����m/G�d8�p��4�`]�ز�?Z��9�h�ʳq���X�1)��9v�G�VPË�hRf�#u����F���aM�4��B��*�a��FX���O� !���짹<����7��2�i8�ȡ�
$�PnT�.��e��y"}_�[Ȑ�ީtL�SG=�o�9k��'�B�ͮ̌�^��Uԝ�Q�����r�Y���3�`�� ���B	������q$F�y�$)Kw�+ށ<.�<HӏB}�%G��'� �U�G}+�fL�D*�m�#�˝y�a�[���*�^����/����x�Ϟl�ϏӉ��ٜjqn2��8�]�N�R��*.[��o\p�� X�@ݑXe=��7��G�������_*���r6�b�&u�w�rO�� ��jR��ލ����/y���"M�w���[`�W�`&�kDI�����ؒ/��ݐø��I��d	vBe=�b����Z ]���<�ϑ�� m�{��趶���N���z�����>G&�l�]5�UcV�wvT�c��1�������`�U7ί�}2kJv�����]��9���-2�-��7Q�C\X$�bS췓��+|�xv�nI��kL�LQ"r�E(����|,H��&����܅�%O�L��;��oz6�ej�`�G#ż�wz��b=��\ĴC~�h޶a`c�� Z�y��l�vr�t����Vd�tF)����I���_m/H)f ���c%��K'NL�W`*�����R��y�^4N�b )����J�V�Et�ܕ!�C?��*����J�q�c�B¿��6'�鞡P��T���/�����1��pG�|;IL&4���l��i�JJ�M���|���A�0t~��:kZ�Іߒ~���]%҄������R�?>>�x��&�L��2w�* �_�(��@�[�eʴ�"�ЅTdU���'n/�x��Y@�q�P�/��'F�9;�u�ӿ�
f=�۶�b�y�Ĳ녽 ���a�$�����j�Ko���|�������� ���[J碼F�:�h�.&�H5�~�I]�S6+?߹<K��C.;hoP���?��U8y���#��;�7$��ǿC��w�d9������7�m!��[��L��g�L�O"���V��`5M�l�	ZNƳ��'ި��ڵ518]WB�=�B��h_]X3ޛkR�3/�&3U5)��S��w����B�d���FJ;N�{,�,1S�l �� >4qEa�gm�`�׺��� ĭ�L-3��R�@�)+bκ[hpnB�����H�����z1��ņ���8E��;��h�x:n�l�ߠe�d�@�^��������/
�S{t��������U]@jN���e�qVr�$\9���T�ް0���Q%<2�_\d��;k�(s�c-^�jޒ���:�B���yt'?�T�&�r�Q�0��˟��ݦ�v䎊�AI���N�Χ�Dk�  �O�/�蓠�hO�3���	dƂf4�l�
C�)=BZ�$�<

|ԧтd��t�D��bXW8�X+��K^��E�)����A )w��O@!��}�<�҄�Lv�)����W�D������KAM ��Z���ǚ���T�!��x	�*���������';��깩i�Yvd��r薨��-��m\b��P��(�!��i��ȕ�)|��f���������i=��ֲ��u�un.�aB3>vԼw���и�,Y�N0�5�x��V'��=�K��=�pa�|pfE�@w��n�^~��,ྡƖ�$�}��,�k�6��dJ8��oMG?}
<�㓫5G�w����0Q�\�A��'@�6Ǫ�t�H=V+��ޞ�W9�>њ�%k��(iu����I��ԯs�:w.�������v������Σ��Cy8¬$M��w���͋��d<��x���}4�
's��/���
��ظM�{A�c���d���#`j�N�q�)���4�Fw��n]�Mz�(�I�"0�����mW���8��y�/5�w��DP:y���.9����z�4��p�%���2��X՜+a�]V��-�V{ ���]ɛ�b������G(�́��n�w2he���,�yXH*�9u��e����[�S�
�"e��:RA;t�ۚ)�"�Z���j���G5�H}#�	JP�lv�+��)@�O �s P�(�"��s0�Q����� �����$�h�Ѫ�O�K�F�j�1�xS�d��B��azM`�"����{C��+��)���7�i�:��5�F^�����+B_�8oKT�x��ǜ��}�GS��.�_@6�֭�c��P��o	LJ�
B<�O��W�)6�=���H\jC���C�F1y"��32Yz��*۵� {.n�\�+5繏��6�zE�/-��2�'�C�Bp��ӥ�8������[Oflc����±u���2�Ǔ�L�<�y���e�+�q\�&��J��������4OON&@�2��P�Fs�&����kⰃNk~ݮ[�'@��%D�nWW̉�b�	�����`���X�Qw!p��8:�%�s���,�;���u��`�}AMx���uo�`�2�{���ޫsw��G��CY<�D�@�WH��x[���$^�.��	 �3T���q�b��%�0(��)�	m���>d�!�1�I�1�LF'�T��Qw�%Z���	T,wS��#��3�� �s����5�p�jb��o��0��|F�5Rbg�F*�<�T�����=VUWD�j`�7�;�Ƨ�軹j�7x2=��X��딝
ᩄ���M�wb4*ր2^��Mz�jX'�vC���,�X'��h-�E��Ay� ���� "a����u�k��׆V�']�g4=} m��`zbOW��k��C ��GeU�2���%�� �`�����ܵ��l��F�j����������ZN���BZ��a�\�)��������@&�Z�h2FΌ���nk�H�p�_�������ƵQ����-��Fx��a�݄���˿�6ڏ�h�w�~x�Q��ڮ��E�&B}��FoCĨ��*7���N����"�d��r.Q���j<]���4����=���!,��*s\�����$KU��U����AkMw�����8>n�=�!�T���0�;�&rg�+M���!���UrGB�k\D��k~MM��҆� ��`���H%��>W�ǵ<�by@Gs�.6e>�-���O[����4
����Qb��x�ш&�N���iy2����\,���Q��Nɦ:A��8��%��_�>��E,�#7�Rݓ}�3��3
��nW����TB���īO��+k,��\D,Mӽ��O��
0�(ʑ�,�w�4(�q�B�����ϧx&@��ͱȀGd���4�vYd,r��4����=�&3ZC{D�r�g)��B�������y�GM���'M�min����M�0����	�����G-f��,�Ǘ3X?N&˙AU��&Ӯ��n�)���I�D]_1T��J8���X^F��C�4�~�������YC����<�*A!Ree�f�F��?�{:��;�_hE֡`�>VW�����EVa%X�����7��!���l� B�����|
l]~�X���\/JGT@,�4q�BS+4$�i�!l7}C:ѣ��?�'�L�Dk}����\\9݌��8.�سM�/t����5��]u�gm�]L$�F<�(�5�M����� W�	&ںb�R�U��nKQ�i��6t,ΰITU��R�R�@��!_�p��k$��v,���������ħK���T���peB�)���dG���eߚƓ�@FnEn]`)�Ƥ]�\��:���R�V���kw���� W�L*��KG4QM@�m��#�5���e��&rHl~a�B~�́> j�~M�����6Bid�@�Q&^J�r�(HӨQ<�ff&dN��X�iB؂�"��]�1�$�w��禰u�0�Z����əZ;�9���(��bǰ��(Rm`�p���?G�O���4���������`��U�a��WuEu��\e��o���Z��>���zJ�M�}y/0�3��
� #,�YH\̴f:7z[I��d;���ӑ�G{tXnC����~f Y�/Kܘ�F~Z=�i0�JO�U�M����u917�g�ǈ���f����?���J�2��6��G� �櫆�}�r�FE�4f��?�;���m� ��Y�j��wdD�' �����]ɣ>F=.-����x�E5O�=��������,��1\�=�C�����I4��P\�Y��8S&��� iũڦh���e��id��)0��s|���
&��M��2�S�D�sCCl�;0�BX�]Ex���Z��_76�8ONt<6��V�;����ðR�{�x	o�nI������;!�L
X��ow�-��q�t�¶vG�����̀�n=4ɋ��]�C#$�/��{�|��->���P�W��)� �[6�U��q�风��E�t�0���˪T4��@MF�U]:���U'�z��],9����8�����:����C�8Ŷz�|��틼v�p�HQ0P*��8Г@Y� ӊ
��#�Y���vm�l��H�u������r��M�Ύ�Ȯ3����Y�ӔT}[�qژp1��n�^��ɚO\&)�,�7?/�MU������)8O(��gM��6����`�a�%�����(���	N�_u���`J��G0�I�f�HkT%�q6G�R�v7��P�#��t��]��^���ȅ��)��L�����"E.s�|(��P�I����yS� �9�{]u�34^�0��_ _  �M�7k��)i�Hf{HD:��jcy�&,_�.��a�c�m��O�{����>w�Q*�F����wss����,�?�w�T�b��\7l�@�òol�������⫅���� �v�7�����(����=�ߣ���>�skx�)o�N�WD�P
L��l5��ɱƯf����U�N����@/��.J�:r"�;S�7�bA -,F.ǿ��v�Z�W���__��Rq�Dj����h�Af2Q��=���Y�&��D����)���X\���?T�ø���7nɴSF��։��~�;���F+�u߅;��p�r���_��K+(�(]����=S�K����g�W��9 �X�~�׮V�C�$8�
l�#r�d9�6�F�Fd�)E�RK&PR`v��߯<z��5������̭�6A���[ǝ��~�_��A$�;�4r�%�̚��p�S��J��k����������H��Eµ�>:�'�0����綧1nC�C'J����Zy�\SB��"FMd�=�R�"� �_�#Pzib��%�lї�>��A������zUV[��5�.�f,9�[W������g.Q�f���n��_rru��=5v���9��uH�/z�|kV�a���RiI�]zv����H��x� RAw���B�K����(`��������x�L��р!���Ch�ູS��*��=9�ɿ#�`�$W�8����D���=�K��,�"�}�GC���,�'�#�a^C��vl<�}�*��-O�ț�~X�u���$�(�=_2�=�����1=��UE:uP�����<�f�Hգ��=W���a�-�=l1���T�
���O�v�/{i��uH%�Y�X�@�R�?NQ���/�H6�jܯ.��?уg�~u<{�[���kߍ���
3۩[{�������4�{�Fu����eM�ٷ����5ӟ]y��]c�n=I|Ը��-������X���+�y5̎�Ì�%�k���4����M��Vk��o �����{��7�{�@�"ՏX�U��4U���٤!`"W�
�Pa�����s�V`��!<7�V�Q��7k��������_O鷓v��?�23C*6",�<Ƚ����q�k��I5	��Wi9�wM������s���c��;�U6 ���a�K��5Ǟ�[k�Bv����+#�t(r��!������8�8�휏��y���P"7SZ��wJ��D�f�b��+���B���3�B���E�5�䵄��O�#��x�o$x5#�X������Q�\���8߲n+a��2�FW� �.+�1[q�iߊ����Q,==�Ju�鋂��m9�]�7L/7�v\Fa��y5�ɛ,��8�!Ο�l�Ćav�&$*?{VG��8�U
�u���C��PLj��S�^8@�{4�+P�8%�U:2���c[?��~��4�^����Z�p�x��l��p8i���/��<тӖ�B�iU�W*R�H��������5 �����A̼b��\\��L�����N	D|�0:*�Y�&v1�^��x5�%t�Ѽ=⣹�6'mT;�>C5���ճ8ӪiS���9� �
���P��?
B����i�ͽ7/=��ADFȫ����D_������͘1�����������b������Q��� ���k�S�S��ó���\f!�t'������cy*��*�r{8I<�4-�#{X���=�p��U����_�-Vergo4]O�<RO�]1���7Pd�Á�3#J��,bLq��2��i�d�4�Yn8hQ[�f�(J9����8��>�R8�U<{lKyg�֝�w6e��)���1�9����"�eʥ��y�����M��ZS�6�+^��L�:�PH�Ig��Q%(eL���t�0�z����k�?,=�#(�mJ�(8�m��Q��`����?�<L � A�a)�rf��g���~W�Q���$I�N�HV�!�UE�?gcZ���A�#ѳ�?F֫Y��ă(U���/��h!�C��P�L�,���VG�b�-m¡.��1�_�z�J*��3U��Ԩ9;r:�}'qga7�k>ϧ��<-�^B���ۉY_��Q0qֱ�	��9��Bi�2X�K�x���x���$`�i�wr"@���*㗺�|�(��)��b��
k6˒�=���bg�3���O�Ҩ��G�B��,���P���p}��":2�,�b��`	}k{0���C��"hI�z��$T��=�m�P�v�4R��-ĈY}�p|H;��ƥ>Le���no�'�E-mk�^�5i��Y0!�ɲ�l�۲�]�pĨe}�ݮ��)��u3�r���3ɉ(�H=�df�il	�.������=��r=/&�q����hɹ�<	�2+:y���zu��@@���1�J1m�;�~4A<w���������<ݽ؃�:A9?��)Ơ����jrMoAH3K�݄����x��|78�ۗ�a��F���z�zHO�TcЙ� �v {(�)π�CؔE�z��I�X�&��ǉ��l���wΓ*���.�M+$�}�� �1�j2�;B\�`
�)���9�WTg&;�C��{X6ʟ6E�����0�9��\�d9�X;�rO�ЖH��fv���|Ņ��t���Pd!��ܤ�����͞W�
�8�󐜔Q��Аr����3۩&���'���9�����X�$'�~�%F/
 ]F&LtR}�W���RV�-������.�U�vQ{�=)�N~c��1p$^U0Un�����<�Yۥ��.'�J�E]~�@t(�m6�_���" `v��A�{%64�N��F���g3��O�B�W-��,SXY�_��xPYk�1��ܑg\��v�F��{�]�*���A�1ׁ���Ip���q�|��W�PH)`O,��`�L/Gx���>�IWdum��.�����R��]"��}�!1L����~��$3MqP�))v� �9�ݓ�g�ʥ����t¾�Q�P��!ܭ�T*�!hEA��0&�6l� ǐK�|\���A�̋u��p�F񛳳i'�}�^�����d�"��Xs�F�y�ȫH[���:C{�v����^�a��:%(��+��x��Ӕa�h��?��K)���`B��e�w���b��{�z)�JҤ�"�r�sdx�%2qLMP��-P�)���f��ޙ pH����/hw��2�l=���,M��`�y�K�G�ݙ���,u.G�^�3X�c��4�V��:c�����OM�������1ó�-��+�+Sg`�@ASA���l��W��8 �.`2���KFTR����BùB��e��mFy���2�a�z�]N2�8H��� U���+#:N|;ν�����B�ne����h�j�|TF�;���D %�t�����Y`ڦ�Za%66'��9�vma*�AQ��sE�4\�*+����>��ԛ��6�c�Q�aw�)�6�Ɵ�z�����8���M�yMG!��%Z�d�g����
]�%0����'q���xU���M�i�ƴ�s��e��~��u�ޖ�%7PKcxC��I���D*Z۝���� 펖�E�_���������)(wō����&	��v# ^)�)I��5�Saq�$��/�.
Bn��PCE˭�k��h��<P�<�!۰n6���V�cK>��앝Nq��1��P��#����n����`g��2L�y���O�Fj���̧kU'����<�{ڹ)UM�&�ȵ�j�'%)k��e�/�V�[����׍�z�����u�{-[^�!@������αQ�r�+O &3�J�H�,�ɳWc&:�.
�3�������P*g���R�����Z��5�<uibM>q�v��ѝޤ�u�'*��I�����(kw ߍqj�n���4u�??�`UZ�i�t2<B��UQ%�����r�(r����׹?������zE�vq�����g��PN����������m홟T�0��_
TY�i�q^B���r�|��±p��p��;5��S3��@e�D�� ^;,���Ǡ��Eʢ_mje"Ҫ����sG���pH�.���P[�|�x����b���X��k�Cv�&?�x6�H۵����r�/��aڈ��Y�
���cS���������!�K� 0=>&�S8�'�q����
*+	���9��@w��xp���
1�aT���Z ���b��l�H���/X���lB�k���{8���&�V ��eT������$|a{�*�#p��݁1I�Ow����%�������ܧ����S�LU�;��fV�O�3��/3��U�?�����H0�Ըv����ʍ�ϩ2d�z� v�X�3�v����m��	+�@���Z��o����0�7�y��[�Eǘ��+]	.�WE�(��x����U���J��_��5$�(P	��i��辟G��Y��<����V.A�0��k��~h~v����bhM`y+�2�"��e59�.��rqw����
�ƴ��B-�5�I�"���%/RK�sԒ�i ,�8l>vD��[ձ�ش�|ȴ��	5/���F�Qp[V�[��X��+��@����9xs�)m��l�b���B�y�9}�e�؁2�*$󘽁F ��~0X'�X����ʘ��#���"D
&�p�z:��|UȻ+�u�p~�%�:\��&���{�upR�aEz���P[ɹ���$aB�i�`�*��*	��b��~y����N� \8[��L0�����+�J�:M錑"��e�,���T��-��MP�q���ɋ�r����FQJ����=�ƀ�&B�Ɠ%���[����:�����9t���+�^6�|�>��-}4��r�;��^�/j�"��G�@�ݮz&�c,,8��q�e�%��70F8>/���
���k4�[��&���'����?��U~y�� ��8RFWtٰ`L�����L[�Du����>��{z?B�0	�^���zM���n8���@J)�:�o'�e��:�&�W|��Q�(��8��r��l���1��g����n��T����i6�r�)��VYh�8<�mϖ���X��fT�]}��/w�����I5��gqG�>{����p�)�Z��Ymȩ�a��)S�nU�j�!a�?�E_m��-,��>���?F仪G+���BVS���&J��|���޷��@QT�~���#>M�[BY;LT1Q:u�߯ǘ���߅�Qݞ��U�$�yKk� ���-.��&m�4cJX����/+�1cS�h@��]^��b��P�C8
�G�E�������[1ZqNef<�_�;ЈCnK�ĀU��ۀ���J�g�$؏E�9�������F����i�0��?�W$5�\�ټ$,q�6'/�hA�P!9�>1�܏�u��]3c�����s��~E{�Q�;L&�����K�%;���}ȅ����mIj�@[K^Œ���e[6Bd����9�aAK��i~�����`���d�t�m�j�Bpae��J��gl��u�N�Ar����0"4T\���o�cWsB~��0F�ѳ�(0��H[_�|��!y}E�T��ddj[���vO�b�p��ɕ2l��Yi��]��]��>���U���v#��������DL����l���^�D.Y�b�
�xm$f�iHw��Ј�c��O�#"���4���aK;��o�A��Px�4J��q�x����[ ��j�)��X��m^�[��"dD���w��,��Q�J�,�-��e�_��
��؆׃�Pk/���~�.��ŕ}�	~�2:������?�gx�A�E�i�؈���cf=)�p	MyT�*�YUÏ���w��Zӯ�<�p(���3�C�@���A%�ϗe�v����h�T[B�:�ҝ�hK��|�����赨V��L����3�(��I'5�c�~�NF\���}�w�Z� 5��dE�L�1�o�e�k��&���*�-���RPN>��$�6�6��+�U�ZX-/y��G�͏X���6��Y��*.)����8fE�<й��I���S[�P�߬��Wq�ZɺI������9͆0��ruqBc��o��s2!]h�6Q�APXIp\	�K/�P|��"��h��x?�.�5��ʥ{"�ÓGTA�i�Y��İ����=����.G4�����x[6�غܠ�l|�Q��-^�'�Rj�"����VFۜ�Z�8<�%j|d����<�'��8��HNY�F��G=�"��>�9YKp����D��t�*�̉�����y�Rl��B��V��"��Xkv�������vyZQ����3��c栠dj��Tpۼy|�ŧ>�f��H�-:��t�qF)ƍ�PZ�[��o ����>ѠE[y��{\�2��|Ar�
���C��?�Qm���l��6�߈t�#t��N��m�"��m��	f�@t� ����w��_�����'Q�� �K�U&x�⥱d����k�nU��g�f�`K0��-����P��W�C�~Ÿ�����<�"nz���x�X��R׳Vb^_䖑вAɟ��xB/���.%ޏ��� ��	��\%�K@�s~��o����(�ݠl�k+מ�g��h�eJ;�^G�`���;n�ٕ�kV�Ӕ�a��ٕ�(��PҔ$!�`ی�~%�;Fb@v�21�׉�)���9�=O�$>�<���������6w*A����rvQ~	�{�pѿ�>?�zT�A�q�N�	S��4�bD�Hh2��4�>�Z�P��n�x߯{f6eyn�q���L�h���$����f� �;�����x
M�~�|�o����c��.�5�_؟�I�,����<�8�iďꅦE�>�Eڨ'mTgiN�_K`�m���K��s�c諟7���H��Nڹv�Xd*�:_��1gn�6Ø%W���M�T���ê�X� ���(�9�^iUSIФ{�e�,�1�:3���lc�;�=�d̃�����0	6�OU*^X�n�I��0<�%ǭ��eR,8�K	�ou40��+�%�Q������G�����o%�,M�ԤPw]�w�h27:5j>��ܯ�j�3�4L�[��}��Բ|��|F�O�Ś|��ŏ>Әy���3�ti��4��\NE�D�bxyw�P��i�|�>V&	|�Y���3�'����uv�PcQR�&��;�k}�Dj�7҉w��*�	H����H���!�!��d}���8#�e�g��1�@�F�`�L�| ��� 4)ދ��	7�u�z2<4�*3���ۍQړ;5�S��[�1
�ڪX� Qmvx�W����\��:b�@��Y��f�~�����y%#��͉>�U�,�d'}�,VH��*��"�>�V$b�؈�,��S=��Qu������8'cQ=�cr�%w:%�i8�t�# ��=0�OBf�f����]&CEFz�m���Y��a��<���k9z�pKh���\һ0Z�4�c�J��axrn��,��S�4���s��>6fRt�I["����2S� P�Q�P��p�{��K�� u*����^QQ�We���a�,�����N���yt����qWF�r�G�Ŏw����sF��y��Y��9�7Zt`Mv.��mߦh3���^��
��?��H퉺K��<IϒI�+��~r`��}����u�9���?1�+Y�����:��Jr^������"1�\*�{�G��)^cv�׃��!�q��9,ue���*pK�6�+9�@P뼏$X��[0�������BO*.�ȄN��[�K�Y�`�0����РE�!��)z Io����I�}l'�_tF)�QD_ӕ"Z%�r�v ���.�ն�bՔ
2�]# �?T�� ��p���D!Ļ��A"uF["@sM�=�8o�t#Zj�0i��s��ߜ��!ai�Ӻ�8Ą��c�]-v� �I�	-����1_gN| �����C�.��p�@]���~>���g���[��|ᰡ-я��%+��.Ip!��L{�{�j,U=��%d�UF@^t-��Ml��#T�Dv*��B�O�,�����=8�/�>9�8���5<n����".٤ت�S���Og���F�r�����M���g-1����γ־�{2Ɛ}��ջ������en���L�k�t���ۃ����b�Dd�3pAN�L<����fX^A�+���%G��y�b0�V�Y�m�+ȥ����^��"om}t�^�U|�ʍt�6Sl����q�kj�e�X�����6��iu���H��Pq&��1!�*i?�����l���m��g�V�Q	�3>�y��e���4��}x��mn��ҧ:��6�vp2A�m�/���"&���tƬ��]q�7!x��?Gm��Ԓ�VFc�!�=��8�0�b՗���@,��2��e�㳦��b0(x�4{q���x�f߲��>�X]/_ *��e@�HW��S����}���Ԅ#:�%�I��nJ3@6�� O�Q*�Y�o�'�LTya��ƾ�����-zrFr�!0��3��F�D�4�" o d�s�Bœ=`��ؠ���tɵg��(���K#�v,.��������rm�V�E�O�)�E
�$ؽx�*OD�!��F�.�N�4Q`G�h����^u�d�	��3��P���K��(�m�����֍䀐5�JЧ�J�� }��W���ep�4%*6R}�Mm�ME�4Hys�ؚ�*�I�@�fq�G�aGޚ�\ |d�ҳ��%�j~dAa����v��Gԫ���eW]F�
��oTc	ya�� ���Yݲ� @�ǨL�=>3�Lg���F���Q�`ٍ��n�{#��+hZ�ڼ��Юpģ�
k3��\$\危�������6�������d ^��W�Y�0eʀ����v��e�Q�~�+%~%	�B���h�}˭f4��%cA#=Y�R̃ٶ�O.�\va�Oe�z6XM�ſTd�����yu>�Z���3t�^F�PUb���-�9�QC>�!�+���fq���W���:�U��Տ�������P�`g�K�������b̝i�����[X��y���tg+ϓ��_�>9����3�^ �ޣْx:
�q���B�>���W�'�/�\��.U-_�Ij����Óu�7b���i��N���t�	��1r��}W@B)��Zt����9��a�Bg��ZI'U�T�p���+�g}-,���1�D�$9����8�-L�����@@VB�B��1��M�,�RU��GoFo�X���8v ����/�%_�������U�UE��Ϸ��~�it^� }y�t� '
k<�Tjʘ��T��e�Ji
�z�e\!�JʲUݔ�R~��(��������*o*��.��B���Å��ͭó|l�=d���ց��o�I�̝�x JV�W��ΠkQ�;��π".A`I�9H��p�ߵ������Ll��T�b��c�����/2�?�qh�G(�- ���hG�
 �����U͖�(�f���?��]H�Qb��aI�ԡ�1���i���=1�p�U&h\.����j��m�EB��>���
���r�A����|��l��)&kqJS��JsQ��4��ۯJ;��Пoۂ��H�7̳�h0L]=��e�M�Z��,�Q|�SC�}�t[����ʳ}��k=���>!V�$d3��@o��DŞؒ��/��R�0�&DĠh�#���u+$D(Z�4������jQk|�w� Z9�'�+8�؂(�������Lt1"�"ڪ�������FX��JvH���w7~��=�q��y�~}�!/z���"~�P��l���<���E� p��^�����.�~�]�����2�{�)�wx�qIx|F��jE,����I�^���4��FSGT���E0��7͜T3kń"r�=�	�SfSxְ� ñ���)���}��"����h���\�z1[��'1���H�F|�O[�����;��j)qz}��*%��M� ��[4�%./N1�@3�<��0���˿�:�^v|#w��zu`����%po��&Y�,���:�F�z����ȗ�ܐf2cA�5C��c�.�T��H�t�Ԓ�κ��O0 H�˯)|�+�9H@(M�AE �Þ=�tp�%1��% ��-��q�]� %c�"~2�]SfWs�1����Rh�9h\���Wh�xqҟH<	�Ͳ(��q]���BKBR&��DZ�V��F>-��q*Ƶ�8��	t��q���U��{�x�n��"�(7���}$�l��j�6*���i�������g3R��YM��Aa������AM[��Ց��&������2���_6
1�wBq@�Y���{��l���ߢ�vxs;w�KԸ4�m��W�F���+R��y�`_�e�1w}D�)��#��.�C^b���u�t��}��6�]�@{@����;�?�*�3Å�!G7ܵ�ew����S��)�Y�j�N�v���2& 
�U4pVWG��ɶӝ1P�i�E�����=X�P�B�)�2Q�
��iD�@�0,�_F*�9�!~8�z��}1su-n'R�+X��q�\�u�\���j��]Cch�=�{+3ƨ�L�{��ȵBk,�C�K��w"E��sHh�'#�J�]�=��Aj3d�C	E^��.�Uu�,p�iΝ#��M���M��9�8f��a��H��vˢv(��[a����`��O�s�b S���L�W�t�z|2��ي5��Ίb
�Z�O]�`p-V�#5-8�?bRm��S)yԊ��
���ל�ƚ.K���{ё���1�ӵl���:ݽo;׀���e�e6��-����4�N�D��7f����9)M����A2��1������U��|ޫ���&I�s4���&<��LJ�R�����]��>����������4PBy�c��F�&�+`�y�p�1�ʂ6�d�������,6���_�v�p�n�c^�^HӚ(��5�,��{-�m�v�v�M+�Y�t�c��l���q��&�@���>���s�R�8���!*���6�6X��
���-g�;&=8�I��|�X�w�F�-����7����!��T9�1Hw��Ζ;���6rz���7�4�+X�ϫ�;��t�[�i��e�_ֲ&V�(�G�Q��@CV��1�'U�p�?���;�=\/�T�x�M��m��F]���S�dr>���E��4E�I�	ޯ#6�Ťx6T�r�7g^d�_Ǚ+�.�#D$���=��.0���M�r�x9"v��h��Y�W���Y�R���z�;��R]���NԠ;|7��H�zۮ�lk�Q�[��=���l��7P�T�r�ԛ��3I��������k٭�nG ����wڗ�F�AX���q�LO�`��>��=�ē�\�!.�z/=8��	�a�a�E��ZO>�������L��ukD����47o�O��|��y*�Ÿw�<�-b��Lp~=���ݷuH�Z~|*�F2#��[ڑ�����"�y��� 	����"��L�oӾW�t�t�Tĵ�\D�7��m��1��:e�#�N�~��O4ھBbӰ�77�%( ���C��P��:��CF=�a~\�8E�w{#����!�؀5a�W��͓��ͨ��`�v�F�
o؏3����ѷ������"&�S� �=O���ݖ�$��ּM�p3q,d��a�c�6*�Dy.u�+�·fI��H�ڊ�B�4+��ۮ,�#���:�0��ҚX�ǣ��`0y���L :Y����@b@i�����}��ds>B�:Sh�L�v�)���Є;H��
�������}�g衴�NMi���ī�9>���LI�=����'������#�#�$kc�;;�'�8`AjQ��އ��K�(0�&'�_=��:D� ;L�I��ofC���wo���b��?_�<�d2��'Z��S��2"�N(��҇T�$�r��)��T�F�qyF@0��.nǣ�Q��y�Q��h�Ռ�3�d?7Z��)K=����34��W�3�\A���}�<¨g�'5ԩ������ 7�H���;<��-@9dx��}|�ѬZ���Iǚ��ڤ���aD�jH澵7��@aC�^�
�	�m.B�p͏s�5��G5;�Fם����A��.'՛�Y�9<xfsn�8��w V�"��Nab�~%]'�W�,!U�>��a�0W�k�>U����ɼ��S��S�����fV���`d��z1�v>� !��b|����H�PU4����^�7Pr�K���������&�=�7,�j�WZ��Տ,S2���مTt���'8�b�q:R�q��4�w�K�����=���0�D�`iF�X�S���aJ>kn�n̥hI�Q�O7��j>Z����򇇵$A̿9a��k��RNk�t���ղk&�kQ�C��ր���ͩ=A�h	�i�������CuK<�:�<莨��l�^WD(X��!k�#�a]c��ۿ�
\���T�������}��yt't>���\`�p��F��(�h���b.Z�=}��GS��B�.$�nǬ3��Bg￡ͥ�N��\L�>��%$��ދ���i=Bei�8�⴨z6�JW=U�����·?��ʲ-|���M��Zd��:d�������8 �e�]�S-	1��?�p��5�ё�Fٮ���(݆}׾���"�
�{*8j�9�\^(�l=�V�-[��� �-�� �� E��.
��ƌ��劤�^�:�ml��o�Q%c��߅S�M"ˉPd|=����Z���@SJ�1&E3�8��w���� ��̀B��ʔu�=4N?�R�$�Yp(�z}������S�����T�wf�X���	�Nz̙�H�r�Xl׮UO^�3գ[�8ht�BJf��ؿ}"���``��C�T�ruz�Nv_1�/��H{o����.�*i_����y�=�rn�o�l�t�I��p\f�&w���Lߕ�b���f9���:D_t��b'�X��dB�굥@�q�f�:)t-5�b��eʱ�BW�����_�e�W�B��v�A�y��k�&Z:/��H�O��Fp�0x�>�ԝ���m��v�U�{[�J��[�����}��H1�q�x��jT\�x����R~���;��NR�����G���A�����Wi>J	�L@U{ {�2�/+מ�8Ux0�*D�+y�oS�@�.�����֮�J SV�q��%��zHX�ܟ��j����l̓ө₮��=����Q@�.����~��]�"{b��J�Jϐc	!�{�IFd��� �f�;D��H���r�����Ѳ�w+$���m9���(�S��w?Y�Z�$�3/5j�D?��nHu`�Gk�_ż�[�Nɨ��a��<�~�9�ޝ7��:�zp�ۛ ��ȧ)n~�=�/H��^Zϕy�����wb01�qx>���xn�#�j�%�4��-�p�{��5n{Yv����
5�:9p_�5"W�h��[����5J$��so5�v��6����
��
��ߔ4�h��|K�U���#w��+�^%Ƽ;��,k[����DFU�kI8��3kL_EkmH�S�B|貺g��*��Զ��@�~}��p��N���{�ʈ=�{'��q�~�=�T��h�/ yy�)c��G$WrQKb,�� /�/�U����M�Z26��oNW��T�U��!�A���	���\p)�TT�g1�1��c��w=$wKwcr<�*�4g�����c�ը89ǘ5A�2�_�,�}�/~  c.������m�q��fe��x�w��LǏ���R�����yXF�U_e�1q&������r���W��V�/�C<�����uz���5;?ؗH���ء��af�Hսfl���y� ���]��oOg�� &_.��aJR�u���Q}�.C�?��[t�Z�Mwt�Sa{|�Mc�$�$=�W�p�	�:�����}e�8^/�4�D�)��;셋�f6�:�k+y?�����x�}�ߝJ[�����{Ȥ��yDu�,�L�t{^B5Me7�dJm���.�k�*:)�V��QAʧ�|�L�6-q�s����'gO�/�%�r��uSceڋ���мE���Z��O�!D�צ�� ����Z�[���"7�Z��6\8H����:6���~��I��$R�_����ݸO��ډ�9���8w��P?�,�Er*�2����f��Z���
�ǀw�n��k�
b�z�<���t�/(А����[��TX���9�א$$A0ѷ)�'X�}�p�n}Ǆ��RR�m1��;Q:��g�:���j#�L�kDֵ�[�j���nǴ��c���r �z���͡�����E����2<���}���;(�z�A�F5��$Ϸb�c��ި+�����n�S�����EVG��p���d,<�}��+վѓeC�r�����M��T�h��� ���HQw�}�3]}h��t�cǶl�����`��R���y�q\�P�&~��6���zs�!��Q�J��ZjC�$rڵ�g�<�(�{��,1���t�)|(�����$Lw�qk{u�]�͠7��-b%�$���J���������@�Q���������A��|Q�<15�>+���d׏��6Cv����������oh��Ӱ��}[��vʣG�F�Ҷ�*�x����Y�����c���V���>G��7���WM���>\'��i���j�O�|�"��>�x�Lff�g@re�ߵ��gQ\U�6�扽97ќ#ghK�s�f*%L$�̒�$.�&�.&��ln�4��Z�߾JkQ�c��HB�a���YE�VV�NIrN��g%��h�A@��b�\u��0J]��k�4����J�&Mz�$\꿓��N10�K�g�7ZWվy�`a���?2�xBϭ,jk.�ąE8T���]1h��ǣ���MY��?���K��l0 �Z�Y��/���t��x��ܟ0/�۱E0#�^�u�mz.�a�G���2��x���Y�,}�F,�$�����U1P���]Ɵ���~A��3��.�ڈm����;3tO.8��5�B�T�2��w쓄C�D��G�vƃ)U��s��wU]?�Bs�`H~uI�zvk���P` ��n��<cA���4`�8̴�r$e;F�Z�f��<z2R��|uA�ѯj�P�,��[�7%N���0�=�H������� ��#�:T�Io~�ۢ9#�"9Dc�:a���f�<X~��6�B�\�����̩�p�i�J=���8K��'м ���a^8F����� J+�Cڃ���C�u�z������D�����٫e�b����ֳ{��"?��C&����\9�I��_��)���[��`} }�g����v�F�F����3߿�D��8Eg/��!��+#��9�b�ɔ���.|CWT����x�@0q�>>#^*u��{�0��t�&�NkR��kqqo�Uل>�?}J�h��zF?.$�!��gp�Î߹��v�oBF���K~0�"sS[T� yϢf��.a���S�����Y��L]���Ϣ�:��dK;G_�F,ۯ�\zX�A���7�qj��qA�
�ju?�I����䄟�ʈ���c��@���D8mE��2ُ�zr��+�p���	S���^�o&��&�xΖɢ Q�ҽ��+�S��2�X�.FMWu��O�|0������jE?_��ez������T��Ө��W'.���	����_�.Kid�z\rB|��.H>�r�Owލ���UW���f��Z5�WQ�A�Nςa*�Kd�u�=��1]��X���^�4ͪ�1	��T�(��)#r!p�/gc��մY����Y��8����3�����t����&<��W����[c�;3>r��?��*<�L���R*��Y���}�,VhrH�ax(�Y���🕸=���-i`�pu�Ҩ�r�l�C���eP.�+n.�6}�h\p���׀ѥi���ӏ.�M��gbp�(G�3��'
)����N!�fM��_�&�vq�K�˽J��C-���^q�2��fa(�{�(A��t��T2WW���I�l�8�Bnya���ӑ%�č?y�lk�
������QE�K6��S���Ɲ3���)%��|��f��$��-���U+��l^�k'�,���U���F�����n ��Ce]_��w������I(��J��(�b��w-	��sBY�(EAwu ���ŭ &�"S�^���?͐��_��E�Ѽ:9�p*�����h_�,C�4�\1\#�-5݅� :��Y���vy/C+@�Bn7�dMq����Mt�w۩��I#�j���X`m�!�1Έ"�RȇUP���EMs��OW�0�=G[~Q4R�lԲ:��љ�V�\K#;ze��>:������g0�Fx�ynl����TGΏ:��25���d���1k׈E��D>Si��8n�~�d���i1��C-�f�T�Eh�`���b�մǉ��ʓx��Y��`��rmT"��0 	Թ:[�����i'h�I9piJd+��G,	��iQ�]Ώ����z0�|���q�4�O���'��F�����8l��@S�u��LK-�x��Ck#��u�T����\M��=��$E���􏈇��8qu�{ᘳ�ʖ��tr���q��� La)� |���;���g3��ʺ���Q`�q�{n@.*|Gz�N=$f��l${�&�N��&��$�⑃Gm�נp!Vh/��O���	n�,���}�s������C̆)�߆�&���S1����k@���Sr��|�cq��X�H�{5�t:��m�-��O�K��te���UT�%=��~d��a�l��y�u7p�E@if}p�k�|���G�4�["V��Y�����
ڎ�U�F��c�$Mʝ�io@�z��ϝ��w�~���-������3j�jΥM���@����H����$qL��_&ff
����6��&�>7�����\~gS����8��ƻ+��{�&4�p����u[��+��M�	�u�F��uE6�&�y� ؆�i֛ ��\�gV�~̐����T�j�5Qi�$,^`v-�-�-�ɤ�7�����	�N��(�O�N_�2:���_�j�W��t�më�ȼ%��K(�G�
Ę�l�:����v�)��t�=X�U��Xȑ���8��o�8��$��YҶ��Wn�xS�:vA�
s.��,zj����e5��HGh�k��Y�1uݮm#���ڋ�h��5�:4��[2�x�,�5��ׅeT������ƒdPF��VCb>�d�[N �4n�"8��P���Oks#%�t��~b3k�R��p�	�9G$�Au.������b��巽>6������A6������k�R�K�.8�Pb�?˳T�`��%�E�E]�䜌 gh+\�����~�Pbtq;k��W����h�NU�'3�E�j��F	� ��1q�\׿��]���%&���Xz;�A!�֟|��d+�V8��@�U=��:^0ݍ ��)d��0*# 悬����g7x&<X���A�L�t�lx�^��W$������:����&'�h�xy⇊��L�{�_×<���g�٬���"��}��x]��/���᝽⺛,܊�TW-��q�<6�u!�����L� �U�,:���U�bŠ��!�ilpm§�p��J�c�ߝ,�YW���V���GL�<^ex*z���U�]:��jb7�V����9�g.[�^��"��[�A���fbZ$��n+�����k�Mb�ۅ��&��f{����y�oZ�r<FՍ�%����׀�[R�\���Ok�JP�&�p]��"�@;Ř�~�4jR��mf�Q/
h�D��{��w��9�J��$��o��EV�Z�a>���e<��3NU�|þ	5��	u���%T� ,����j�)L���w�]v*�r��(;^*s�/��匳���'H�[��6���U4���@Kl\�ef�}�G)���T��@׽�?�vt��ZŊ��99�1�H�s�{�e[�-�x�բ�y�Y�TS�ܷ�P�q�7�Op����U�f�c{H�N�挑�m��T�ŝ��+jg��/[��	�a1i���
aP?f�Y�'�\�*���dkD�g��~�U	�Z�V�x`��.;ŋ���DD�lXm	G6��~]����N2h�/�!�����l��z�U1�.#bf��y�8.\�ݕ-��r�if��.�R&�ǲn�����q�P}�6��U:Vî����a�����F@N�Jv�sd7���g�n�[ff�T�4����[��ω�{��~#	�%Tn��	˛�D�W�0w��HN|8_�C�`�XT��ĆJ
�6�@VU8F$���OX��_T��Ӳ{6�&�4uM1�F:�b�x���J�X�Obv�E��?:��9���x�`%v���!�ͽb>XyJ�W�/:ʽ�鈚���d��UY׈p�T����!@�������N��|=軳T'�f��ޝd
���Z*����`t{�ԧ�{0�$������܁ ���s����k1��l�,2�=�$�J�~L��@���E�1l~X�5"���G�I���[!G<������gu)i���~e���Iŭ耟r:[�|�I!{`�V��*Kn�@�,�t����:�G�y\,���s��e u,w
v$���|�W­�S��^�b�Թ4$E�)?P�k���,M�ؽ3 �����h�#��W�b�(R�b�>L/�����˕
"A��������:�I)�&�be=YT��ϴ�@�s��K���O��P�PCr���ˑe���y�2%�9�|iBPuA���u����BçG�1��˷� $��a��j�L��g�Qc�i�YQ���a�WX������G��8���l/�*u�	ﯤ[�B��ֽ��ڈ��"��T�s�ݳOK��D���kf���m'��_���j����pm��7�q�ڙ)4��ە���]�SQ��$����Ԇ֔8L=�ˌ�4���\���Ц������f=,!�eP	�\���[�����+/�/����`���aǗvɖ�ڴ7�a��TLNQ��`�n:cx��3ۻ�#P�g�t�������Z~W)�$�� b��I��M�-6����fS6��c�w%��)WBCQ]�
��D�����%EX8t��T�6��_�|�A�h��3�^虰�Vzhû���"�8k�����	����Z���H(��J�f�gt�+x��c=L@j�q8`R����8�^��|��jı UMJ�䕡&��b��|T1�1/���]���F!��G����,����b�?�P��f��Icjl�U����p:��E*����PW4^2R��=��0]��-��Y�j�y�_?��^���i}�-U{��[(���*��'�}��0f��A_�SW�ŋ���-�p�q�)i4��4�B�f���R_���ܧ4��:gU��98����]�a�m4�5�6q�w�V�E�F���^�u�����xa9��;��_��B�oMr�rN�D[ڨTh��7��HwS^��`�g��'L{���L��ϋhN®S�q�ud���8��[ �)�ւ�^�n���C�5[�<�P��a��L�jy�^��*�r�����߽����{��I.�y�BF�e��3{�7H(��X#����
_����YM:�a�j��򻏅(�&�M���"��0�Wy~�i�5��c�i߬�$?��[��>C_G��-P���r���X�����C{�.���x�b��U���`�e��oDq�\�Kb:�1n��GX[�j��}'#aQ�C6�;6������YR-a�|��*1�ݶs��b�8�`��ԝ$�4��.`������LY'i UXbX�."���Ed�
�n�S��o棆"g���)������92���ZRQd|uO����a�௸�lc#�~�W��^B������`k)���+5)R���geYz���h��u���Ǭ9֗�}�+i�= 7��$�`�T 8s�8�2�4��2�T�#�*��OA
�����h�a��� ��Ww��;�j��k�n�_|*/<B�L�׸>{v3E��|��(�J�����c'���X���v`6�?>"@B�Y��5|̘����7������EF*�	2V������;7`PH �q�i�<�X�Xl��pLB�LS߸��� �o��`q��i��(�����ȇW��]�"�fg�jF1�P�v��x���JV�tH�4L|&G�}��q.�o
���ώo���4n�k
�]&�k=���vZ�f�~�2%��4|�����0�׫9����lߠ̮�M����}���x�f��:����;�(P3E����Ɲ����1[/�Q1�|�(=Z�5N��q���ů�0��g^Ѣo�HI�V�/I�j��_-�S�O�!�K"�KB�F/�	܁O�_��N�np��"����$`�w���ti��>-�y;] Ɯǆ���>��� �}����;�o" �"Σ=�Z)7�F��/��_j���5�!F�����p���zD�C�];�$V�%]#����d(���U%{�W}P�4�?����d�4*��eQS�e�����M=��=����K�]6l�;w��r��`r�����QB&�n[���c/��^15�]D�rm.l�;����{F�=��[o:�z:\�_ǁf��B+�י�a���ꝩ�(�(ż�Yע�:UU!y�������*[+E�誅5:�X4%�p>�׹��!�:�\����t}M�\�03(�u�-d�2��Im��i,��H��6uC��b��#�W��l#[�Z�f$	�<ۑ��uل���$�H)R@�r� ���I��KdP���F�'�����;c�-���9;N�qd׽�*i�M��u�	$�A3��D��Q��#���H��ϻe�i���4I�PL�蠈��-�1O?�ee�_XG/�~������_ ��͓��#Q&��y�_����LV�xm��X��30�{=�9����-��ɞ�>MH��6w�;��сmԢ�:�M9�l=����23�j����O�\�@��ɘ�x���̻����[;Z��L�E��{�`�w��[�j:��[����Zt�	�;t�m'��Z�a�^(0x�Z<����@�C�k��m�K�����Ƣi��(3�j�lu�6� %%8b��鑣�g�A���&��<�<�L�f1z�ף9VK�X��P�0�(
�O�$��g�r:���oǊf[�QR1:�e_IO�ҵbςe���o�@9����V?~���A�0�� ���2�ǩw<fh�!<��E��愆#�Iu-�nh�>���陣}*e������^{:�|�ǗTnt����xl�V����+�#��cS`�Z�A�0��k\�k���(,��:Cn�Z��y�\v�����q�A3�5�x\�S��g�+��I��y�����N�15�Z�'=��8>#��f�I(^�lQ%9��D�C�7�d��Xo�?���='ee��<b�%�8��?��gt��fwn2�����"�s�������a2c�WN+1Q�w��?邠zeܱ>&���8c�E��;+xX�%c5��^4�iL	��H�M�]�p����x�����Ers߳��.��hu�1b���*!�p������n����P��^%�}g�{SO��?��Ui�:�W�T��������_r�0&Ol6N}ȍ;����h��/��I�8\��u�+���
�(;�	�F��#<Dy�����6f{hhvj��,''L����
�Gs���-A��]�p��.�f!?G}s~$��38#ް暩a����������_���Km�ء��k/���@�ޘVd_-8��ذa�'�f�t��V�/w�iFЋ:��j:$��S$�&��ڵ����^�@@q���D�S�F@��lA���- z2�����h�P��#�i%�t�y">㸭YWL��w3o�ՉH<N�[#�� �����7_A���c��]�G�n&)$�x����t��f��M��r2%���BڍHn����KЗ��CGZ~$��p�+�r��ߖ.7r����Ru�)�}5]����֔|��ꡇ�׸�+���Ă�Lei/�\�;���&x��cwJ���_�����,�*�C��А�M�>7Sc��<j����oGD���q�����kÉ��[��z�4�sm��5*m��Y��Б�$��?wa���5�T�n9��t��k��t�j�\3�DͶ�O���V�e��H���R�L���zJ��
�	�`U�1�y�PǢ��E#r���f�pݚ�C=r�ި����1�ՔY�K ����, KW�X�CqQ���Tubj�����>����`�D�~�p�Ep�F�SJ���Tkax�o�a�z��+�.��m�Rx�ȗ��i�xzO�S�Y�z���S�JD:-r�� �7�ҡ��=�j��H���w<�����ѳ_�ǐM�--�0a��Hm�K��=RzX�����h���o߅>�q���zn�����7j�7�]"p܌��4�Bh��8�m�afZ�{mo_qC���j�_V�
�ޙ�p|mX!�C�	е�з�1�p�洗*�HEU7�EY\�j���� w|v�,`�W+7EUC�-�F��/tV�$W�մR67�V_�̍��y�߄�L)0�mC%�*'o��*s�5A�2��'�j��L:�$��6,�~��=�ݬ��-.�z�'5�g� I�?�f��Ű����X��Ժ��dc�(NI;��I��a��Qw�,���CS.� &�:�ǖ�ٍ����6Nx����3`|k�o`���!x�g�odh�8mn�?���P���	����O`���C~j_`�O��u��{S_���"U��D��X!`T�����b@�}�;%u�"v#��Rtn�kY(��BTS��z�e:�!�d� ����\9�V*A3MV_�Z�����k��QhT�ܽ$�v�ᦷ���[�=.�	@-JN����"�X��lKE��8t��عL';z�x�P\�-Z�+�9翬���m+����(w�ڵ��"J/�+e*'��� D��K���I�:Gj���<�⯨B0Ok'Y����_��i�J�#,N��iO�b�w��[&XyN^C�V2�M�����Z��gK^	��9�f듵�ީ���Fc)q�c�G/�?;��k��^��\z ����ܺ��8�ܢ&��=|Jў7�h{S���X
��o-C��É1U B���h���خ�{�k�q.r��XA��m�y._�~�h*���3E|^���Z}oQ8q�FM�7V)|& ���!^�k�p2����EI_���) t�����5��0c�W�9;��Lu��*X{�#c�����"�ʳ�:a�غ�U�k��qvx�`d�E� ��燳+��C�]�����<c,-�������o?bf��Ԁq��M�C�
�GE��ӒF�V�j�h��9��q[�9���o~��f�^�Mc�Ѱ9����bE�5�N�ɑ:��$6���	$�Q���Nk��K�e��B��F�C�V	Ī�U];��w^1��a�)ͪ����Ԇ*�O�P�z�9{�sG[r����
�=~ؕH���::znM્Id�dt����Y�V�H�nb�Bq��9�M;��j���'�jI���Sm/�������gi{�"�0�$��&�K�ш]�X�^�	����b3���D��W"3$Xiz���Rgj�x�O��xC��D>�sįV�. ���oe?�+g1oF�+�˚F�tڎ�qH�U��.@��ߪ���V���j��z����io@�%,u�|�����1�#����7w�MV�/�q���/G���A�[��F}���R=@fj9"P"S�+��̐ K���yW�nhM<�	�'�N��M����Bpn����Ǌ��ya|�+�	�{8j bZp��J)xMĵ 6ל^@�[[`�����-gܔ,��w���v��EF���p��t���l)f�w��zF�H-#*f�C"�V-��(,;0�
G�,9=�2*��l�#�c?U� Om�����T��$�%������98��E��D+ �[���)��י���X�T��Nw"H�5��t�0_[�P G�;4�pd���E������X���^���eofn&�R�}�^���!v��������O?7���@\w"P��-ߘ/��
4Wr��[raH5��n� #��6�!R=�T��zP���y��oր�v�	af&@��*d���	�Ra��+����n���c�O�� X8"�����[����y�t��Ll0k7�԰���\OI� I���^S'ֈ�iX�7j�����j�`�#˷"��� *H�c.�8�;�E��w��mb��);�`.��55�ސOr(ۜg����9VC3�8���<��zb�AO ���'GW)���T$�q\�Qzl�M�rO��fymH�
#Q����j��/�LBS�ƍ����y��ʦ�="& (���Cb�>K[mDx���f+�$�������{����7�O�t�U)Y��Q���_@�yL���W˲��.���U a��+��p���{����M�>�5wy,�D`��d�w�L�GA�̙�I�M��X���Ό��E�f9�XD鷦��T2@B?­��?��W���x[V� �����d�����0	ks�C4O�dc��3� ��|?I-g~��2v���i�#�(�����I�ַW��!���f��|��{p�Ru���ah?�����p")��s�ތ6\M�������Il��\j/�cߩ�T�׻���<��E���s �+ƋLʀ�ZClܚOj�Gԍ��C� �l��N�ɡ�[�F�.m���ҽ���4_��s�0��x�9V����n�[�������Q9���W~du�+��''����f��.��������r|E 02�i�ƈ��iAY������,���42O���>wYaCҊ ���JTڏβwW;��&�w�F�|��t)[6�Q�u&�Tҟ:��y�o�����r���={$05�;^i�F[C��3<F���]��S������Ў��g��"��ڑ1[	�`���[
��r^W> w�JI)a����^t��݂/�=y���z��}0��Z����ֺ%�M�`cY�Eg]��*��������w��o����̈x�8�p���XE��}�N�I[$�jv���D}�tx�Ž�mfJ#�K1���k5���R/����:�@CVR�{Xe�%���ӑ�x���kոH|�JH��`|����;e���r�}MY���ϛR�A��l�c��ȓo<�� _J�����4��m�q��l��7�p�)Gڡ���C�^�_�����U�ZBi�:�H�@U����"��ix�^􋪹o�C@T�֛A�C�N�t���S͌́o@�o@�A�t�
%u��~G ��g=`"Jq�ǘ�VA5�-�(�"�����2bX�\�a���ͱ,<�*��(�����T�
������Н�;3���?/�]�C��oPSV/��6��iE6hO�p���@�3���-xp��v+ة�c\��/sWBi!g�a�$����ѣD�H�iBi����a�3��\3�fV[5H�8�/��[xMh*�Ї:��X+@�4�I��3R��Y�lJ�h�(�#,~ ��D;�����cO�"�+�W��[q2p��Z�{$��~d(B�̜U���$��U��3X�c�ta:��Wa��~KKf��]�V�2�7���A�|(.%!Zs�k�?�h.������skv:�����<T
����[�cܕ��_�q�R���2x6Rv�#���mQ�D�K�R����c���Kn��҃�Ϲ�j�F�,θ��6R����U��F�t���m!�Ht-���0��͍���w0]�h��e��N	l�Z����e~�)D��gE�EpB�����20�B}z���qI�dk����j��/"u>Ϝ*��,����a�j�� ��|̲�r[�����0�Wl(�{�#l�u�s�U	T� �������lU���P�������A��Y�j��LؐNQ�qO�b�߫2���*�}�����bȀN �M�D\(�R��U-s���Xc�eY�kT�T�}�q���5>����(�Mg��U˸03�1U<���1���cr5=����,[4k�E�]���9�ʠt�Ij��^V�t�_��k�(�FF��������kܭ ��[��T���+FV8+��r	J3G����Ժ�_��kz��1�qm�2�������c!x�
�|"��8�����SUyk�Z�m	"�ZǼkr�:Yd6�F��a޺�)�C҃���A��@�g�22�%�2bR������2ޥ�w�|��S{M���
i2�����¿o��N��r�kפ��kՉ�V���]�|��������U�~���3��O��S����� ���yǆ�j��lm٠
 .U�#Y l]3�_�_w�zNf ν�����Q���P�A��K�D�+oONj@V��� ��ս�j�h��OqΩ��&L=�|"o*�1�;"�-����o �v�fg��P,cm�|�<|� s"�`����z�c�|�Ac�<�>Xv��)����4�SI��v=p���:�*�?��x��*���OV����I���.N�!0��� ��fS��$,:f�-��%n�Y��I%PE�^|�n�6�[�o�����4�߯�%��5������R�i�*[\0�r���\%���+�8M�@ ���Q�yo}�v�{�C~��#�� ���DXP" �F���KȚ�~^&�#񣇮��	u�Q�qJ����
݊����U�I�k�O�_z�C��wP��c4�6�eHT��jp�_��	P>�R1�T�?�9�!�I��ol3�r��l�J�;��Xzi�Ń�u��ׁ�x\�'�>$�e̵�b��x�T�N�gMڡy[��ؐ����x����hG����)Q�-�WX綫�6Zձ�p9ҝ���7� R�>z���S�jb̈́ʟ8{�}F�a����e�P>C}��$_�;���gOޜG<��̘�s��M޹�)�)3%�G�P�(%�1�2I�6B&�8b]EE��r~��VB��4�V�N�.K��_a >APRp��:�����֡�yG�4��F�^E��R#k�L9[���0zoh���NJ��w�FX��ۦ(���%�����D�3��h����^��M��Ds�$1r�R]�;��kE�ߥ�'
1��yb��MZ�_�:�o�_� �U�#鶬���zC�a6e�a�E0�N���Y�H��D�&y���!>������oÕ��p�n�X�[)M��K�շ��y���e��np4�����K��2m���F�� �uv?g�k ŕ����r�������9X�z�kwwi�8iash��͕P��q,�s�)?�H/����*�R���xk��x���}�|"b��������b����W������#� �u�Ž�ǫaG◇%�2�l�(UڪQr�P\'3���nK���S�M���������Aq�5�"m[�=�*V�eg��r(J���R<�r[��b\���6K���=@�JN<�I�(��i1�9���a$�g`O��Q�d�چ6"��J��6�~�����@߳2��(s�n�ن��f-��p�[4Lb����jA�)���|:&W��J�}�rk���Ó��QM�l�vIᡶ��E�ё��t�s1pr��c�$S������Tރ���#Z6�?�����.�@�F�$$���4:�g�2��D��0@�����5�c0E�_���u�k7=8)�܍?�w�5P�	lw�{D�F	!�;�f ҕ�2�+�8[���X/�K��6�s�XL#A��PP3�V��Z��V�)"C���� �xΘ��׈|<r?l��l�6�Z.��m9�'��WkL �qd��)e�8�vw^�Ɛ�b!.��/��c�Q��$6���������׮n�_zh�(�b�$r�b�ڭIh3.��V��Q�e�B�2���g�{b�Ud�c��SH.%��ŸVla�C Q����R�gCE�?-��l�ʣ� P�Z���d��H��o���*�<��� �����>�X~�0��V����[R-_1����KG�;��}��r�CBZ�Z�4lp��'����J�{��I��,�&p�&4��u:����ы+�S	o����J04�����ٰ�9�fjP��8��#AH�����o�9�@�6a�ً}�]�(�ga Bc�w7��<M�!�	�$� A�QхQ��%PY9�J1\����0vn�Od��S��,�C�mN�_U>���Ԏ��	F��m*�s-�^�2:36-�~1:��D�C!�]\��N-9z*@�<,-j���9����e�7,lx*�>�K�d�,3�t�V��KoX*$'�f��4[A_��B�^���W��-SȈ����,�)�a��'&�hT%`'P����r�a7�5��hUS�:h�fh�ϫ-�析 �JSI�TfQ.S��.�\L��(3A�E�&���W����u�I!R���_M�q+�ŧ���SS,�u�nU�͇����E�0_j *	:��h醹k������F�d1�m��>!���v�eR�x�p������~���o� �pn�@��3�_��e8�Ҧ$�VSR�P�(�J12i;���.y~�yvζy�{�c���p_M#��dy���"�ǣ���������a���A��� ++�_IF���`3��c2<x'�_�x��AwI�	�~���Ժ�rXox�e�e/N=Z�LV��n'���1r�I�ؿ�-B���t��Q�%j0�2���@R7���.xDK�*�)A�d��\%�uF;��H���4I+Gc�^��;0b�=ծ�h���ϩ&��
��X���C�UL���*9&p����&�e]�K��m޹ד���0��ޚ�����b���{!׺�ro�yИ�T»b����gȡ��;�P��4�����9�,=	߽�&~����B��_�7{Mb+�R�� �3)-#v�!��q��)2={L�A����7*�=W�F��Ξ���#����fp�4]�P���Ո �DҦ�ܯ�q5�S�E��~��1�����j�M5�{��)��������2�n�,?�i�u ��HRp[���Ӥȉ8�+�0o����p�w��2q(ޝkQ��w� ���?�*�A��w�f C��+��v��YV�[1je�p寳W�����_=�N�����Az3t
�7U�۴��W�5 ��U���3����E$��C�� ��}s�u)�Y�xp��'{RĀ7z,�U����҇]�����f
p�,�\M���)�n�m��[�n����m	�ː� ��6X}x�㿏�]y^��皛��F���ɬ�d�"�:�5D�4�)��ah�׫�k��_�X��\S�P~�Ԝ�ө�o
]��\�[�� I���>�!��~$K>n*) 6�]�h<?f����4I$8$����4%�@�)c���}�sֺ`$[�n<�V���)�ʜ�h��y�A,�WV<�|��Iz"��/�(�=g>�}�f�g�S
ur����B�'�#�|r���:M���X���p�f�7j_��n�0�n��G�v L���Lأ ���k˭��Q_+ڙZ;:bnx΢��և��5M]�m������b��b�o�i�~׼�������I&���q������|�������5�lv�9­�a�]��̽ܛ �Glp���5ְ����z��r�g1u�'G]�hc8��6��}��
P��|��nFE9��W�fh/��H�s5MR����(Sԓ�K�3;���1�!Dǌc1�S����o`h�\�Y.�n��-��;G��1�!�9������Ѵ�i�.�ç
O�٥����w��N�c/)b��?"S!tO�Z�®������h#M���n�R�Ѷ�(c��ŝT�+睒�mz�-N�fQ�;Ò�N$��� �Ez�u+��;�#9�l*�L+A�J�'(���H��f�<�ǢG6C�����F[�ªs�u��\&��TWb([���0?y�!�#B��7l��B"n�\^��D���L�H���m0����X\�� �'M̳���y��ُKK�z��o� ���ջ�0�i�Ҥ\BnY�N��nQW�py[�E����&��� � ��:j��rdo���<�^�H�����]L�U� �-��د�.�+dT�w���	_^���� 2�_A`nΖ������g����|��k��L�v��ܛ+���VN-.�75S���ǦY����yٟ�͌��/��������,�V�v����S�P����;`B��G�Q5��O�g�8KW��j�!}���.7����H��#*j>"�X+!祦�B��R �s0�e&��(ey����c��������2E���T/��ٙ�mK�d ws٨�:i%��{(��,��L���T�X_�z/�q�?K EƁ�o��e{������\SAZ�6;A?�#u���S�X�o��+��IvZ���%.����甕��84�y��QG+����R�E�l*��]�>��Ɣ0/�8����]?��Bb�ĺ����^���=�mGCP������w	�,�a�� r�|?�og�
wľ����м2n(fx�
6N�Nݚ;I'#*\Q�<o���K���	-��>����{�G�n�f�2XW�e�G�L��[û���:-���H`?�YA����~��-D�B�P˅U��U4m~�i���������y8� ��|r��+���,�P���p��u���>�BUZ�����h��7��.��,X�S����'��p]���@{g`�[nB��=��.�M����*-Ox/�� V�Z��G�p�xR�t�vA�ֶ\
�e\*���!d���8��?�T#�S�1�;J���'�^���w9�[̗�̗�Y�Ȥ�q��j���b�!�v4��A@M(���$��E��]�B��{��q�s�ߐ�<������	I�Ƽ��i�UÆl�>_I��jٜEh��i ]s����t�J�̞R��A\2���N��#�!{�kxg1�p���w�ta?�]<�:/_����Ll�K���*�� xz,��-d$Q|�"|�VFﵟ��n�-Z�PƐ�^����`+5��|���K�=�:7���#�J���D!�v"�3�U�jj$Ԕb�?Ů�^j^��x���dK����	�=�]�]ҵ�4:�j>%��$��'�Eb�c �q~6�g��\��s֙��Z��Y "��L�{�!�oN�����9�3��$K�S��g�&��+.�b V���e.�%o�4������a�#����P�`�kt������T�dC����񰕮xJ6��4�
_��ඕ鰟4�@����`#d?N�!��N��n�F������e����T:D���O�:�T���,ޑ����J����1!t�ߩǒ��5���K���L�6Z���V$�:���U���#,A�P ��~m���8�GM�X7:����J�`�����ܝs�� �{��)BWb�v�:�2?���o+�{�L,C���0�����o�rsݼ���hD�@Q F���a�H*������_��A���t�ˮBʊjy�؀�[?�o���?j.�KL����4����%�_�N�������ն����*R�F�;]ܼ�պu0�
 ���D����WY�G�y�5�5�7Th��]~�>���m���G��zVxiRt%�� �҈ֆsR�:yk�A��n�'�J6W���{c<�M��o�6��z.�8���}Zz�C��.bC����~�6g�\��i�*� �V�R�(��v
1� �'�@/�w�x�+H�2Qvr-a�}�RXE�'�A��pC�gF}�\���}����&I�3%	f�=�KDz@d��L�J�r(�8o�w���$�	�
�:��s�=|{8���t�D�y���i��"P���\�J
%�>D�
�UF����7��.��e�xn����0o�e�JAZ'Ɨ����!+��)�E�D{�͢����K{i��
�ɼ��i	Y��ǃz1�*7�0N�u)!&+�:T�nSKhU��>)nEğ�)}#��B�� �;eM��v��ۂy��l��g$����o<Yee�A�K�~Q������7%��Ȋ�󫨠�����{%XH�8P&��R��
��3=�A��N	�'t�X)�1H@Bׁ��+g���a9�~���LWx�F�R�˕�� �b���㍂��5�/~��6����#.��"d��|�3O�Fm� � �+U5Lϕ�=�"��'^�ES���E����3	6�`�0�tP�+��2�`>&=��S]phI�[B*qi�.�@���i��Gh�tb��Kbbe�ۆ.��R>�8e%���H����sGJ��z�L���,�E��ê4���+���"�9 Ի�6g�O�X�2lC��8ӂy����딲�ݺ���B	�h�m��h�b��
�q�����*����h�9;�3�H��]Y�#6zJ'd
�����e���+=Bp����,j�[q93��#������820��/q�f��i�U�� �8�P�JuZ'�&���E����)�{������v��W��Ăx�O��*���rD��D̻��H��ti��O�j�o�{!)z��Y�zO��"�bI�Wx��u�2�>E�ҐK�E�
Dj�+K�	 �cW/����i�q�����{�"�0	���OC�%bG1A����G��$�hh�ͧ�9��k*z�w�D��5�`f텷���m�D��G˩��'H�)�#��xiS�AHt](W��̇:�z�l����o2������~�g�j3��^5=S�������N���k �dt%��.�?T��p/ހ)j_T߆�����mŹJ��T��{ʴP�H٨	{V����O$��dP�F*%��X�c3�#����&T�^<<w���>B�<B;B��^��0!� �T���~��2v�")��}�����~���`�'�3�0�gD���(���s�L���l��T�g3�.T%�����\,H��	��;� Qf�f �
i(o<�f��@�l�-�&�Wt��JD� �Y���ڔ����C�j��d���"�BzQi(��O"�o�Yq�%�ck���:�J�Ne7{<'�=m��)���=�u�A���md+�`	��l� %������u���ϊ}�"���Lm��LB_�Q��,�'ߦ'�G*�Ŀ�D7@PWɟz��쿦8�Y����dp"�yI���º�s�l�q�VO�Y[p7��U��dR�H�k!���Nk���}�WK3
-��($�Lݕ�>.�@�&�[,��V�I�h�i?oބYD(����/��MEy��W�M�_�<j�!�����B�s���sWŊ�G���&�ߐ�^MbdSW��IQi��q�&�ia��1���D�T/pQ�n���[Z���j?�w�6uۜ��Wg��?��WM	OA��V�Ux��I=j�&���s�H���Q���G��>(��|�^��;��)$.��:��d�:�s�14��i�����HP x -I��<��_��Ϧ����	������̀��'�Ui�b-Jտ�R�
v�*A�;���Z�&�j;�{te?��V�#CZT1��n����&-�%:��������~��!���߈��ds1��w����1v�Y����R�}z����%d���0�`�`3�-s3��V����[s;ń�����f`8fm(<�n�4�}��ȱ�-�i��s �y��h��@�]��&b��L53��k�	�2�J�9�����&�o�P�JFC���@�BL���_؍�¢_*DV#v��Tq[SZR�Ab��/G��m>HJ��~�a������n�U�o|�����N�[�&��I�L�ug�q��B��ɸ|�)�#`��R���3����1���X��pf�Ϛ#��"4��o�q��u��n��V����_-J�f�j�φ���rv-H�P�<�kg��l8~��q��y�xu���'���1p���x���2�K�'f=e7�M���~ʩO�f��;U\<n9)I��2�ŷ)���`,O==ck7�)QpB���
���`U1h��.l4;��i(����?:^�Ga�(xOX���F�B����+�CM@ę��=d��7f}�m�E�Vxx+�΢=a#
�w w�gI2%	s���l?��Pc�Yx�+n���!���������SO�U��i��K�Ő����J���]�h&�T(ʦo�R�3Qf�D&P{n�Z����--��$Y�J}����B5nfզ���@���qA��П9�Z���t�G�	iW���\�j8n��t�������0�X��y��<֤rH�R�S��#��DE�3�j	�u�#t�܅�r3��U��a�
�n��P��2M�������2Gct��"V��F]:�-��>[��8���Ud�� �$};W�
��Y�ڢ"����ץ�� hƔ�{*�I�z	0W��_)��i1�
F;7�6�
�(��y�?��&<L��lTr/��3`�N6Uǧ���n���>�.�^K����c3��	d�����W�~�����D����i�0����L?��=���hX�"��S���/nu��Y�B.��03\�ً�pt��P-� �6�VF��{���J���O;�'YB�1bv9=�'}�E
�
�c��дh	����aHL`߸jw�G臹 8�]�tw �	�W`���ޅNg{�DOP�37ط@�~�Y�*��mI��+�N�&a߀���HB�A���d��z�N�����"Fs��1؎�*�$�	�rۓnv8(^���F��nZ���)��`FG�|���&���8��4N�Z΀1�nHΜ����(�Q���ƾķK��0ݘ�f_�PhW�������K��À��<�g��|���+]]ނW޷4|�ۜH_��`�>�����`g
�T�9����tz�
�zg���yрG��C�e2%�v�pD\]5u^�^�2��6���Q�$
ZY`M��Ks�&��8�}���uqu{�)b �\Y7�CrTM�[�[1z�������_����g�.� ��_ojGk?�ʊp��j���	����Œ����"w�|9;�ʘ�b��uD-<���P���y3���fo�(����	�c�zBD�)��ϓle-᧲ �d/ډ�Ǳ����(��6ׇ��`�;k:8񻥪f7{���i�έm�I�z�l��^�C���	_{��a�'��A;0v�8���B���p���3�SC���� �B,�p:6 �Aq�MM��7��/�4�U��+�i�0x�X_�h܅��(Ƃi��?��.��9�z�F�\�"��������T�(��岫BtlŁ�Cn�y)��q�r�4�[��[��&>�b��3��ݿU�Dl�!�V�@����+��Iz���ǫ�+�*�O�J���+NyTS{��R����ե	�$�Z�ͺD��z:Ȩ��s�h]�y[��<}�y=6����� t+��
���A�j�u�0W)����^��z"hpWBvT{�w�!�]�j��%�.��f��?���u�s�Q_)c?�Տ�n�dl���L2�o-���Y��^w5E��Ï��9��B*�$R���	,�;�:m��i�#��U�xhB1��M��hhfŇ:Ih{{�l��yN9�H���jDT��^�+���&"�^��HJ[� ]�.�@��������H�ý�~��z���=�.x�L�AjX��W�3�V�����g�����/���۪��e	&c�:����>�>��K*(>up ����r:*��?��Հ�y$ױ��i�@�˭N�`d��J�;*(����8O<���Q?\[O�c%Έ�"^tT���ǥ =J���8����! �H��A	L{-�{fc��:Y�G|�5
�W3������ֺ�;�l0�Z�l�m!�T�Z��A�Yv�9��M�=}�rC��H+�b�_
�����)sIk� � 0O:C��0�I,t��!�I7eoTėɏ��i)�F�u����s���X�梉�_���fI0}����|���'مRI����wh�Zٰ�)������$�܆��ki�1C�fΨ+�	<�M��hЂ�^\��~��<�»3xBǵkźV~�[��I1z1��ȷU���YM?��"�,��`c�<���-82������gfC5��W���.�5p�[D�������C�i`t))B��!>�T�'z���0ML�u[���j��_�#A����M�*���r�U_P��RFE��=՗��6��$��8�ؐ�����N���k鯾[��
�y{�J|���
���束���J��U���|�f7j��:�M��w�4\O*�i�1�^r3n;=3-��2�e��^L�I���E��*��ܷ2��߷AV��	�9����hd>]�n�n�9�鰠y���V\2�TX=3�@���[2
��P�<^�F����]��5��MKK��cNX`�6Gk�4�i����4����n�}4F�����hH��|��kV�{?+6V�� ����<$�"��>�e+��s 1ۋʿP�/��(�������h����{l�q��G=/�Xv�˨x�R=���e8Iz�-��{�~sf���V�ܕEj��(-�q�"�˃\��rl�jY%t���~��e�>n���x@��j6٣�O�VZ"]Wg�}����!��n�>b���QqvJ�7&�X��7EЛ=-9�>W鷓�E=k�CS�p��s���57B�K���7>�L�ȭX�E�)ƍo�}�1K�M�Y�\����c�飤�u�_V}&:�*w�:19ԛRM	�r95e�q�a9B��z�$HG��!y8�����}�ȃs`�Z6ik�a�=-����X*������q8�w��r)?���23g����Q�hFZ6>��&|Sk�)�^R���#���A�&!g�A
	�ElPs~-G�b['�����e�/y�j�-IL�w3��
W��@��
(}��&�q�ZD��V��"��]ꡖ�u_��Q��\� mƂ�&�{���u�#����'���W�v�v"�?	���}�?u+ ���،Y�H6,)Y�-������6�+��l�'�濅��w�<TV�I|u��Kb���ĺ��;=��Զ�����L���Q̐� �
����L���\ǥ#�R�hQfU�p�,�����H��J�z)�_�Sz ���nܰ�.|�RBw�Ra�X��r���vd1,�gu!J ��W9�
��Gж��mr��Eo�6_G��ma��bD;Es��~�v��f�@��Ϫ��j2�����5i�|SU|�6�D%ȃ7v.�j)�`w�)^W��s�?��g%�gvh�H�&_�3�\�]�����IN���� o�e/�8M�_�p�g��0�3�h|PcX���b;K���V*izW��>��˱���,z�s���7[R��-(��Kmh���k	�d'1���t�?&a"�4��6B�姐3'M�Z`.[�f�Gr���=f�.tGmQ�4P- Z�r��T�����n��n�$ ����f�X��/��H��j^���}�'�Ot�O���%Xd��&��~�q6_R�KRbt*��0��uO�{�Dq<�ǳ2)���Ο���)�U�98P��eE,�hC�J�\�4˂�::a���+�����J��<ns���@X�JS��f�ٱ<��q���D1�� ��sR�(O�/�� m�h�Zh���s��VnǬ�/}�95�Q�Сtj��pã��\�L
Ǒe���]���.;�\��ے���`M[N���a��x�kKߔ8wZ����zb��u�*���yj�@�`3l���3e_���݁LXeu Rq�Aa(����^�~�&���XAɚy�-�|%NaSHO7�[�2\�ȅ�4�� �ùK�5>���2���e���a�1-���䭫���m1�c� �|��!�F�~��x�Qlf����탘DUշk��� ;�n�MP����8Er����J���\�o8��ی�Y�����$>B+kI���4���wL��R��`���	����h@¾7�U��v�.'W��1�H�}��0����+�K(5b�҄ʉmͬ�늝��pd�juHV����CϘOj�s���\�6`c��B����������cU������3�l�*�����O�*[��U�W�`��L���J��<0~K�[�IQ�f�XF�s�e�ba̿���Fm���r��#��r�<F+��չEK	�n�E����<U���
�Z�Ȃ��Q��� M�1�/��M����'Y� +vPzM�Q-W⺙	5��������D��'�r���ge�I�f��L���Ɩ�b2��w�Ai�X�$��N�͞	�P��FĽ�?��-p6ы�\8	#A��Y�B@�����י4-��M�h�rǈ��C�^�]c5_�K����dl�3kY�}f�f��>���7�r��ͧ���1��<�5vፁ�s�eqˤ$��mY���YE^�i߷\���/X�a�S�ڄi&G�~�(����d*�1)a�-	��I��b�{��AכU}�,��2�N&m���ճ>�fE��	5X�X!��-#�g=�����B�_]�V��ͥ�� vZ��O�̛c@Ջ���i3�v��j��CG��b�{����lA�f`���0�/����E��Zwb�
j���Wa�r��1�� ޳L��eҨ���\Ef�ߦ�p��"�ٻ�T�dX��UyB �G�.d�FI����&��UO�X�7�m^:�5"��Z�A}�o�$���\;;���1�v=��b9T֐k���·��'9����p�1j�Qmw'�=7�T�n�5x
�����xA�%�"rYo���Gac�῏����{ PRH�l`���4���U�-���mi�^D����&AC)%���Ӫ�*�d�|8��YPcw�,��%����ס|��q�h��d#�&#;���9��yH���l��͛�N/Y�+���� e��S��P>�	B�A�YE�=ET��1��?�e��AV�30n34�i�ݡ4�����d[6��}�Q�ʃQGւ	�܃0�z���]Y(�%�#�/�ETǪo��;�0\~y�|@Lcetܝ� �^B.ݡ�8��cv��KH��Rw̭��.M�XD�N�~��=�9&/�8��8,F���V�s脃/�+��[�U�E���|�1�?�y�gpy�.B	���b�w�tC�).�^�ҳ����2������x�w�漇@�k��(�><�qQn�ǆ}S��WN≏]�0�w��-���\i͈�Մu8 ���!Ր��$r��>����շ,�Z���n1k���+�����Y�!�V���`�ae�6�%��W�N��C[U_LV�#�S���s��N�q�Ӂ��V�R�sO$�z���;���Z"ev�����J��/Z&lp�R�'�~���꯺��["�l��Ҟ!@w��Ⱦƚ�if��+�l�PS���޿��&�[�J��a���X���qu�X�CI]ui.3&�0�%��?#��mcN�PzZ�[:;��b��H6:C<=���j�$�e(��_�L�j���W^Z�~E��T5;�^�z������uMBjF��+�5D�-��{%YY�Zq�E��	I�?���KD$s2v<��Q�i�O�����g�@��S��%n*n��)�'ϵaZ �hg>e���e������F���½����z��?��eѾ>)Wظu�)��ao��:��蒈_��:o�3�e���+I���+�Bҽ�o.s}�HW�~���m�l��J��R?��ޭϤ�>�ۿ������9�͂�ҭg�6���Q%��k�t�n�PA��A��3ÐФ"=���c��x ��$����5x�c�����w��i����,��v��{��>y�S��ONl� f(6w�FbY�rߎ9� ��[.����J�����5��3@��iG��}-ox̯�F\��ڇ���4P�E;�´ذ�枹<q&5�=o#�@4�Bz��n����?��D����8�k(Tӿ0�*��(~�zB��mC�]��ǒ������!���������nw.[�93�Ay�/�SQF|�������f��4	�e�O�{�v����KCIl�
�&��^�_	ᖏ��$��]�O%;O�:6_vP��6�6�� ֮�U�tJ%�54Z@�@�F�v�����v��1���%�DӖ7饷��4�C��1��B4H�+;C��O�1ՒsN@�~�A5�<�i5S��<H��������c�_(�-9�&���G�s��/G�q8��T:s�8�[]��m�k�'I��!�G�Bw�5�Ҳ��V�/HV���1��W��]���r4Jsj%5lE��`�,��}��4�q"�K�xQX�]�X�1�1�`������O�)��p:��j�x��tY�����Z��I�>�Iܟ0!M�A�c �Z��.aa�C�pvnr�)1�%��ye�q`ͥ�T�mFII ���]`�e�o�٪������g8M!����R܉Js���[&{d0 ^�Y�YG�+�h���Be���i�/�+��7�?�|G�-[���g&�oU��&B�������}7^^��nW$`���(<n���I:r���+�uw]e��4r�ݷ�Z��m�D�W�/��I�G�3�t@Ϭ�݊��Wì�m�F3�EOüK��5>�ڰJ��m�Qms9g�Ҍ�)���}��k��|O�Xz��j�J+�X�WO)��ϿG����cn=CŞ�8hs����XP.���X��,�;���z��{Z��qG|r��9��2!���6 �;^�j�S��H'�G(Z�PB�K�������品�`!�h��TGGW]7iy�kTzx$yt��凁Ф��+�Di��b�x^���9]�k�Ȋ��	��o"�i��7�8��d;� .�!�L8�����4T��&r�`��Ύ�n#�R�}]����،��͐v������R�]�=�>H ���'G=�
��0�cfQ1>g��LkQ ��{��-�?��s��/o��W��LS6�f:羍1��T�U��dz�D2WK	��n�y'	��*v�{���і�(@�)o���߽�ɪ�+Ne�����j
��M���}�����bcL��V�~r5M����,m(b� =@���N��ʠQh�z��F!1U�c`N�Z�5��4���E�n�n)ߤ��by��*���/6X�3ًq�r���Y=�T�8�&��EL�1��}�4�!�)�ʦ�'����=���3�����S����9��2�u��@�jk�a�Q��6E��f����JO3E�,�0')B�ٱ��)N��{t����ܰ�6s�@
!l��!D�k[�*M:M�dY��������w3;=�xI���=��U��p3��&��\��HVQ%9�߅��B_��ލ��O 
�٫�����*$�c�q�<%���X�k։��#D<��1�[?��O�=6��1�G��7�H����紥�r�`Y����Vo��'b�q��m��1�-�77a l��Ei�9������ܤx[P�w�T',����[����S'�UB�����i�-��C�+�ݻ��h��4�3�S����"j�\|yS���\�1�!��XB����M��N%)�g2"5�`i�f�������i��O�4���)-7׵�J��!��Ѱ$�(���Þ�����6;�	>�BB�;_;%�z�ZP����w�&��Bo���������1Z���=���.D���$�����V���-�t���<�&����_���Npz�e|��� Ni����V1
@��n~���N�N���9�U��٘E��s�J�E
����sj�)���7�K��a�ҙ̬@�8����ʙu������֪r�c}�����9ܗ�@7���~SS�k�-A9�X:5M+S���Ϸ�ѯa a}o���Dz���7�WU�)����"D=�p���rB�BaY3����f��wO�`Bu
~��m��t+r�7)�ھm�"QXV���d��@��d����+���$�4�Z�?�f��K�Hs��>�wr��
�Pi��a���XC�����xOΊ��C���uU��	��{]SS�9Z7}��S�m�^��,[t5_ݿ�� ���U���6���,��y���Ҩ ����[J��j˹$�6}૯�ds�+��j�|�D����J�۠���I�Yَ��X磗��vFehZ]Ǫ�~��%����4F�C�"fX��+ql�fc=�?DӅ�sF�f�H����X�L���2�3aǮ�)q���2�+�o^���d+�RX���r������Sx��� ��qL�q�<�Vl3A���V#�W����kj�6��Z֤X;:s�e���	�t>�X�c7�g�}���.�H�i��%Y`�� ��0xr��XH�`�E�W�C#�84cg�	���~��X�ُ�� ���q��4�/xb���,�8"�HG��������L���/g�M0�`h�ϸ�C�s�_L&�G}����=\柩0̻b)�����"��	��?����#���	�����7���X�O�� ��������̵A�拵o�Q�-MV?)I��0<!�?��^(?Q������:�Q���̥�P7��S|� ��'uf�A��Ay%��&���҈>��Z�� �y��'XzG=ԑ���|m+�ɆH6k1]���W�c��Sb�tu� @9$|�N�qm&:.NX.�9-��A�o�F{�kΝ���-�:��O�m�UX��.�#��-V�f�e�a��jX�Jù ���s�C%@YS��t�����M�� ���:�/2�aɈ���3�)��h�vWQ�߰n�}K�%���`a�m'�%a����+��AC�';	��k�s`��q��J��!���#��y3��ԥř�ʾJ^3[}�˜��r(o��$��ZɅ��E�(���䔀6삉Ӱ���m=z[�u�*B*�p1i�5�M�����u���4ۣ�-�e�2tqK�nQ6Nw��?����G:�4�^0��|����"��"d��Zf�Ph	�8���8ݪ��o��Էz�+?QKC���^�͖�m���D?Y�E��d�t������DH�/�m+��h�Ҷ�n�)m�G6$�����R(����[͎$��0�C�#���g]S����]�O���X�vqKE$q3s��"��>��n�}9�~4y�B��v��1^26�;�&�'�~!H{+%��l�"jR�*����p:�<��0�-pPH`�,�aP����[��!����S�D��@ؤ�F���Vv����֩z&*�X�Ka=er}�L���ύ���`r�9B��K�ӈ�*�и��6�ذ�_���Z�*=�v�M���nk7Kr�x�SZ#�2�rW�o�V2�0 gڡ��� #o���ͩ��]��J��H������ޣ� f.k��
�raŕ�Ѡ0�I�M~/n���[�����ąì�U�����X�d��K�a�{#᛭`]�c+��r���$��yQu�e�����o4qZ=�z�H�PGK�3�~V����	 >�cM��u?�6!���&`�S�����ڦ���U��q.��>����#�^���4���̬р9m.bFf�T8@w�5��f�����N�v/�H1�$K�����&����-�L�؞�`�#���n�����K��b`�n�6:��f��� /#��"�kKH{F\���C�m�7>���ߌ�3E"��]=�v�)B4솬^9]�~.էx���~1��N�T�捓�5V����H�z�vw��#-q#:����o��ZU4�S�ՠK �����(;H�uM��б7��ή������#?�W:`��h��wy��������<~	JOI\^���1W��/D�����4��I�uE3�	���"O���n���0Gi�.�<�o��,�4��̺`��md��u M}$�9W+/��Z����6�����U��`�Aw�M�3�����ĘY҈�ե�:�ٯ�ӯ��Ƕ�I�d7+���A�)�e=M���;���!���k�&��k��䳖��F��]��'v�V�,.α��^�W�����]��P��*����q��l裨HL��mO� �l�ߴ��_U{�Foa�4�]��R�HI�[[�ֽ�Zt��dlx�c>�k-�2��X_��!��7�1�_�t�=�1���α�Q=���-�d<!�zZ2�`r�{���t�J��q"�5/Q�Xo�H��4�$������6��˹��Æ�g�`He4*%�u��l�w|��ha	�2�+��M�P	�Q�_�g��1��k�h�u�_D��^�l�k������=qe� uȜ�����r�߁��,��2�Q�FR�{o-�[��z^~��^ �9Qx�+�{(<��;d��E��U�O�Da�B��.�w��|���k�Q	�`��h V�;-ˋ�����J�SO�-w�����U���\}�$v�*Qd5���9�`���%�%/ej�,��\�_xSғ��0�H���0���S��t�T @J�I7MF����K�Qy< ���^%����7֑;�oI��f����ٻ��H��_�+����n�U>��������Ȓ�a��pP��(���4�qny��gGGc;1� e�y��]��{w�q�(��U���a�f�|��E���͠J�B����Oíl#��-<�sa�������_�A�PP)��œH�����|jb>��Ý#l8�sHBS1	���s&�cc�t�o#��)�YL�*1/Qf�����~Х?�9��<Y��Fԅ)mP��i
�s��
��ct�[�bK�[�K? xe�Ve��F4�1��rk�V�y�u\۾�Ji�!&_W��l;�iZ���L�mX:�7S9���f~G�jz|/��gf����'�ݶE;uZ{�ٽ��rL�_�i�r	8�nj��Cb��,v���L7��B�ʤ}��ni��!�ɸ:�Ծ��"��럋n0���u=,��Ύb��>u��G�Qt����++MGolR?�4xac��xz����L�����:W��"_����k��H˦��}ބ�K���AȔ�$;�2�?vx�Dd�9K�l�ԕ�z$�&	�]a��Y�(��R�`��$
-7�n<�7��"��:w(<�2;Pj_Ԋ�C$��PI�d�# b�����$d.V�qF4�{�:$�N��?��&��[f/}�s:	�&�K��E	��@b��EAig��$ud
�e��x���@�?��jj �8ho�XX���<Eᇹ�_��x��K"�AIN�Cf�!�|[���<��V� �ץ��
���ގ��颼t��2�WX���+0��q!dK<�'pvp��gxtR\�'�����	�Z�"#.�&���=�.P�Q��}[ְ" ������f�z>1=��f�.�	���ݎu����y�g�q���Q> ;�\aa
܍�Q��^�w^���7��\�,U���)�3YYC�g+:Ϟ�\��5fn�iSAkĻ��l���n�f���b�����l�n�ĦX4��It�Q�2ɗU�$�c*��������Z��@H�'K�ߐ�EM7�I�,?��_I�I�gu�u�ͦ�����a�ژ&.�RIR�%u��v�3GN���x��Ϥ`'~7��b ƙ�u҅����C(T�F�/�Y2��I��ay�c*��ޟw A���Wsq�i��6�X�f+Ԯ�%e��j����-�u�P�:�����;��)�@}�*[ww��� �\����za���l�*;\�U���Ea�x(L&x�g�
�'�����+�CA`F���s|ä�:HÉ�*Y�5���5�z"�au�Z�o =_L���Z+�(Lq*�
��% �q�Xr�����x�R(+���j��B]<�ҕz�8�g�+9M��dUҍ<�4��[2
��Hv�6�Y�ۼm@HZհX.-�7�i�$}z�Peal���ꂌ���'eKy�JjE�gL��<2���[|h�x����������"���_]7XX{�P��9��e�úW)IH�2l�4�? �˃`e�'�2!���e�-��o9�Jd��t�>(|�>{��I@�4_kY�i�'��`��A"���2/�+X)��t�m�P,+˝�l��f�<�,���t�5&ִk�n5�t[��f���;?C|Dڨ=L��l��q�e�[�L}e���+p��6
ߡ�td,�
�c D��,G���O�e�G�r(���r�>�:Xl�`j:�@�3��Ǿ%��1Q��Bg�n\�A�5ϑ+�B�_���aO������,��#�������|$���Co����NH%$&��=2��>�w��"YΕM�����F]���C+�������Vw��� B'<�z��~��h1�^z7s6fTH	b������[>i�.A�"�"�T�w��͓әH�cV�&}�O�n�M�:��X��I�:��$�����*��@ˑYt�P���=CJ�~s-~�c.�Ң��*=�bL�]�C�"���@2~yj<��5&MuR��{ɞ��:.j�E�IM�x3rv�!��x��Ŧ22e�{�ޮFj)M_���}6�-�ʍ��OƄ�yJs<�8�BP��̃.|y���@W��\U{^FNYݩ��p>f��O�
_�A���4���D��F't/������>�n�!��,G$N7�
��3��G�g_�BpW�c��嶏E�<��ŕ�W�`�W�M��Cω�9d 5��bĩ_L�w�iH�F�+���t_h�|�ظM��/NN]�&�����گ	)ن�c7q"ަH��1�.�'B^s$���_�\���J����e._R�"��&r�6-�R�EW�7��,tՑ�}^��@����F/�#���W �r��D��XR6�K�9�OP���R7���*(�E���3QU+R�}�5���E`�,d � ]�����a��r���[;�Ԟ��X?��w2�$C�Y$�'G�,��+��S���*���f�"�)�%j�Φd�[uҟm���$;i�_��I���/ǞC�}�k,S�8�@���]R�>@��K�	����1�|lZX��Y���^��
�xD�r"���%m�T����}
kL1�e 
d�9�����
���o��)�!��o׮s�0ʂU���A�&���MF�U������.�b�bh)c�O{��Ï*Γ��߶���״��X�0�v&��"�	����v
$m�B����������ec���@/����_��K�ԑ���-<gŉM�&n>��T@�R�Q�P��_JfO{�4g���{uW޺�� ���r�2��;{/p�J�
B���P��yP�rJ()WzS�8K�U�V�>�;1�KՕb38�G��`��4L�K;z��zγAqN�'j�Ƒ�aoڲSc�ד��}b��O�s���g�r�#�K��U�y޹#���w���X�R�`ȼ���Y��>����`
�ׯ�qÛ����2���]/�t��"�٣=�\���r���$t�°����
d*~X�y���CF�S�'��?��Ө���rf�F��Re��FD���9q����)!L�x��4� �,0~�T�B㒔�X����3����:[�ės�.[�uT�kє^r�`�:��X�F�A����Yt�Cp����Nv0�C��y����%c�] b7�x�ӳ�g��y�##��O��Ӽ>,7��LCA��a,����A	~~�f�nL0+��'�_��,n��-_��ڀ��Y���sF�P���d�k�ڎ���������������]�=�ؔN�h��㶙��n���{��T�:˘�1`)6$`k0+������\`���Ӑ���< ���_���&�b~�l_������9M�sp�\\+�M!0��ȇ0T?ԗ?�q
w*���|vj�����^���8��+<��לU���yiN����Kˡ\A���A:��c�i�j��t��]�`	0��/N ���<9`\L�����P�8�C�{��f���S(�`�����f|�-�w��_��Yǣ���2y]$+����1fGw��gϨ�Rc؂9iM�y�H�a�r� ۀ�#�HN�/L.F \bL �Dc�e�����0#p�,yq��g{+��J��$�19��{�ĺ�hQi�+K�m�.�k��sH|l����֟ yn��Z_�C��w���~ސ�8��-�?��r�E?�! M��xQ8Xz�7��B���������;�_<$N������$l��W�
N�Qƹ��5V��X8]�{C��P-R��,ma�d�9C�5A� �ͺ��T>������ wm����.#��P�-�'�����v���q�A�wi	GZ68t�����j(�D�云_�\���r``%��3�T-1��	KB2�}>L�J圂��4m�]T�]�s���y��H���i�H7�"8��8@q���g�X� ]��ݞl�/�I:k�֠J�_0D�Os*�▝�j"�  ��^+60�W��*-D����8�M��1��&��>������#���{̆� �\E��G՘��M��"��O�O'�J�/.���/oҿ����,��4�P��A�v����ݩW���5�f��9����Aq.�`=xX�tm���'6 m�4b��0�6�٘l����\\�:]���qu{=�?�|����u����9�n�!h�%��:2!y
n3��Ө���^�9s>�h�ū5���Ԟ+M��
�M=�4�Ru�����~���z�՗r�h/�&��߬���OT���Z�<�
�����N��$pM���{�)e.�WLܝ�+��綎��,�s��d�j�,�N��̌���"����׹��#��㟹����3�G{�>��.V=$�W +&�M�����M�)w�b�s<p:G�Gh�c��W�~izk50��zv�ɺH��$�M�I>]N�AO��&��Jzк9ᜏ���`3������m���H�������Gh���әfHx���x�����a@��9�^����������iE�����8,�}H]f�;�(�$��B-
�����#�Q��M=u	����3p�����9p������� ۺ���aW( ���\���w���\�]4i2RS���Q;�U� �^%3���oǽ+��ʅ�TS��1>V�������`��Xg-�4���U0��U��S�}(_���^��c�@f}��y\�3��Y�"��!�xh���|���
�;�$q�E+Y����:&���� �>�����ks8B.�A�����|_�i/T���'u1�7�b�e����oЄ`WhD(�d~b�͏m��()�bo�~li�DƘ�c�П-A��JC� $�!�g"P������aR`C��m�8{R(�A��ڎ S��?kt����i�G��f�G�ȏGP��c��̞5��8�`�3s����cn%S�j��w���#�"ܦ]	��OL��?�A��F��0ß^���^ӒH&ЬN'���K,)3�6a��c����,�4PVZ5�"��bE���0��?��3뗽�/��|Ǎ�NNw[<��|�a���
���uT� �J򱨎h�I��}j�Dl\�Y�לy.V^*��z�W[��JS�6P�7հ��\{��Zic����T������B�k�A�E��Y<%􉟜kd���m�h����7������HU�Ș����/_֔�K��k��\Ʉ����G����m�|�R��0O��	���	�)�,[yr8�h���*}�\΍�'hf�����^Ta���Xۡza�\U_<��68	�Kt�S2��]DC�ޚ���!�E����G�XI��'��j4�L䱶g��C,B1tq#���T����5�{��Υ���vn��#��+����>x����pr�:(x������(��Ö�y�!�r_5��1���<���-Q�,QonP�3c@�H�4>���1&8�t�"�oS��{O��J/A˭^�Su���O��&�4�J�bP=.����o>@�
������,o=O��|�!�"G[W���������!6R	~�Y*C���
]��q�Ak.���:z:T�>-e�e쩦$��>As�RKP��e)�gzj�ͷB��`c���_S��(�auq���r\(��7�pD�j ��Ȃ�ʷ�$����^�TMHK=�7�$�Q"(�&��7��=U���_%�6U4{�'����6�Rs��e訅��Ym>F�GgP���a~wd�;(�er�T��Y�}��p_z<)�
�����7Ȫ/��HE���e�3�~<��Ϥ��N��e����@_��g�d/�(Q�ѕ^'��d y�E����cE��?��FC5p%�����QԱ��f�#ގ��_�1�F���o���K\(y�R�T0AE�^�\�|8������
�oF/�7[��%�|�w^b�̾�̼��G}�/��O<����:��$�^���!yk`1�fq�_��n��@�=�����g�V��}�Y�s���墅��.6�H�r@��$tm��N�襡��Fm]y^.TK�;�T6�t&�gÉա��
m���*}t53��w�"}F^+�ȗ��~?S�$��$!�W���j�؝G�^�$��g!��i5�R��U�o�rv-TfW������ntD����5>�9�:�iSZ��7>ϖV�2�c�I����DC&s������,�AM�$�$�ُ��`4&;�x3[!�n�]*ޟ�/E�PF�e~��(�U�xÓ���nHM�H�C{Qtt�B ��6������W�
�������#�7���p_�.0��ӱ��x4����_�ߑ:�o�O��-�7�R�>��A�(��=T��}�Rҫ)�gvV���Q���h����R�V7u�Y!���d�����\n�ƊмQ�-~!�#�W�������N�L��T�jc%�a��bt�O�Q�l�U�r����F���-ܸ�B����k�I��}�M�����r�E��;B����^uϱc$��>)o64�c��(���2��Ĭ�*p��_��3[qN��{�/��%p'��I_ KH��K�̽7�������#��@GDh�����@���	O�2����>�;���@qi=���N�J�y�xx��L��Z��YR����>����+vH����Q� �����j
[�8 �;��څ�\�j���-��F�^�2�(�}ĒM�VSu��I�ཟ� ��Tp��T�Q{�=BUѾ��f�G����G��ش�h9�5$��Xy��V�M]��OfظQ������}�mp���	����ʱQ~�F[: �_<Qfp}�&י�<��W��K�{;�ks�pH�3��8� �S�$�����CaZp	ܫQ�%G��k=�2a�ծ"�8���xT����d���>yB`�t��d4�$&�2^ֻ�5�4e%{�:�����[K�.H�IǏrR8��K�� � ���� ���������i�� �x�Ay�ښ��w6�*y��*�)�i+$����7���5)ai�����'Lf�˙zj��g���c�>�5/��Р�r9����;���c}�tE�VPtv�A0��߉��=�+"��	��1���95ȫ��DMsџ"�wh�ˬE�L��z$��/mG�b'\,��սV|DZ���p����^G2���f�xO½�>-��F�Hk���)#1�.��s�{q��Aq߻o�IԊ ��a�l���J�_�4�B����J�>��ʘ���%��g���=��c��ί�s?n˲E�H��a�ߛO��+:�ч��\Z��B{H�f4�y���ǈ�/dH���Ȼ�Gt,����D̾�s���eY0t�Ѐ+6�ؔ0��˞�$���H��J-;�shY�PYؔ�p�����wG��-���T�uw?Vg���'��rM�͘p��UN0���u�Jr�Ҽ���@)��MK�ˮ]<�	D^�Ju��hf���@6N#Y9)�uy'�	���iTw�a����`i�Al�/�?�j{n	��:�,c�A�h��/	2T�ɫKA^*��K�Ҡ�| ���~;MK?�v��s�r��n/ 9��GQ
��W���S�K������o��}�i�\f�0#s"�/��k�x<��`A>�AZ�rx��W�N!�!z��t>a_ߝ�K�'�&P�K!�S��7�)'���p�c��|��MK�b�����D�@"
;��Uݿ0]�GQ���vi��e�/h�}\Hb*=N2�}��k�-�$��ք�*y/�ZZos�4R䟰D<K��ߗ5���Н��^*$��oqY<��b:	��{�MrO�����8iR��U�^迏�%0�!׭;sa��ER�$"RR�7��_X�h���t�~	��ׂK2hFyK��9���E�d��ӓM�ct������A�<��}�bk�)��;�V���8hd-X���J�ҥ���?��ӌ	� +�{�/g���C��`�֯,��A�T�w�>�򉋅��5��\e��cbӢqe���<C/��8���r��2�GXCr̄��N&Zo�p�K��ZH�����#'��`wtin����/$�{��q��*/v��A��]x�������	�������b}Hh����˄�
�B�rF�"!��]�4�J��(��-����	��h�g�?ɌEö�CE��p y����3F�U�]���E�A�l�d��*F�7�N���c� ��[`����r����-5��cԿ�,�; �κ�<��O$̜��@�gM��h��z(�'��B4Pp�έ�� ����!�\O�e��6޴烿���B�l�����T���{ے�5o��a�'|`�������&���O�Ce�~��ko���S��I��-2J
5��<Z7S��b鼧XU���/�Hy6A�(O�rI��0q�|��ug�Ǭ�P/�u,��6s%_����VԆ>ʹsw�f�X���N&|�)4�^Kԑ�uPpʤa(P�����%@L �U�� �9N��/�m��߭��ֻ�^1G+��]�'��,� 1���O����P���s��[�@���	��ָv8�ư�mm�J��#�h��s	|�f�_�]��-X�޶7\e�O��u~�P�!����k����f�Z�lg
�|�+�ImrX�-p�(⳨��C�&�?g���}R�7�7_NM"�z���6ԋ��ѝĜ��^jiu(Za9�heK ������)s��=J뷑���C�ltF�D���\�a:�L��gN���*.�0�4"C7���,E�G���"���D���x�9�7I��.����ي�v�fy75G?�ר�Y^u<k�(<�B�T��rvL�i�;�[�N�H����O�]�����U�Z1N/�^��ȆΣ�*C2�m)ں��ׅ�i��Suw�����DA	�	Y�pK�7;*��P�X��a����q�u����
�ń�)t���g�x�������(R}�#�_{������f"�8U�!�K�dŦ"H���*�`5��D�t+�#|EQ�~Y$��������D���_����|��앣�c���)X���<ֱ��ZU�J��H�v���mt|GM=ms��x��t���j��Nʦ�������<���D�O$s����<\O���8n�0*�E�	/��x�|���<$Y���XA/�᭫����s��텪���a�Ճ?쇣ߧa,�v	�j�yw�6~I���N�Bu�ԧ���Gp�����w�}�+�$�A� �>�lً��Z%a��?��36f7P|�Y��ş���1L��b�Y��B0J�ViF��S��.\U�3#���&��׀R�vh�7�s�Js[�xq $,�3PEA��Mk`ߢH�U����O����䅶�?L�<�V�/�����M�.�|����v�~)�k��N�
7�ۺU�x�#��'�Kq��S�$�������'yC7S�6�{ϖ�����$oK��"�V���M�p��֚�6yV�\R��L�� xP��a}Q骮��K��-FA�<^^1ܹ�k.C���E�,CR*���f'Ь�&�u�;2n����E�G���d�#jI�e��{�~o�����i���f&�`
9��^x	��׽��yBځZ��#gȚ������F[�p�����M!����ɠ�w?�?�tXܷW[�b��i v2ػ�,nC�JH
!���4Hr������O���O���7��� nxFb隔��X�>�=�q�۹}��g(c��0����D�7F���+x���U�5�?4�mȑb��!���z%?Q��
\ƪ*�ٟ�C2p)��^M�/���Q��'�3�ms�����#_�����aJ �툨����p��bc�h@�M
��m�-� �գ�={��_#��7`uw���]O@!�OAQh<�ck��t~�B��W$�,���By�n]��w�wrɴ94a���'F�Ar�J�g�cR5�J�fڙ7��%i�!P�)��fޘ���5ǴU׺��כ
�T�zSQW1:�p�Ӈ߲$�A۝��Rfֽs���`8#k. ��p#N�u���U��z��uMy;Z&���EFeF��F7���.d��⃄<��9��2�ӕ��cA�.4����&����.ǕޏϜ�"����*�M��Uj�<v>�� �	0h2�5aY>5a���{7����y�p�a�[�Fd%�oͩ��ᩤޟ�o a?��:��W �� �����Ϫ��m�Is��<j�P��3�"DX���������R�5�}}>V��"�g�	&���<���xt�����T�!&��pࠠ�s�jY�y����cb҇�������.�v�͞�N�B׶���J�:��$�
��T]�@i4�5'�����q]i�Ѩ��"��⍋P���%@fΞD[��Ia) ��ܼH3�]���^4&��f��mn��T�X;�w᫈*��o
3&|.<{�̐�wk�U�R*$��i�'���Ԛ�a�F:w�l�å֔+�?^����_�3%c]�J�qز����(��x�kؖp��c��[5<�q�Ė����H���~y5�/�a%{�"��WC��5AWn�-�,cr���x��6cU#u��ߵ�+�7�u�z�༥��ߔ̙���C�5)сǒ� *��g�k�gP�p�vfFb�7z�^���E�.��\w?".�N[2�?OǸ��R��wS���4��'�=6y(�8��+	���!�WС ,�����>�	��@�Z��lI��ݞ@Z��H�ܽdY�Dl��ϟG�a�E�o�2�a�Z;H�9<l�(�]��b����¦)��kCZH�	�����|�Tօ��d%\�
�-���\x�>BSZ����{Pڨ~*�Gk�;4��Lр|��=
�to~ g8{ĄS�����P�y%C�����>S�	�$���\��6K?�I63���	"��:Vj.�;Sa;�W�*$)�v����L��<��yX0��	i���^���i&l<z�0�a�?0B���.ܜ�+�N�h����.3�����r~�qv�qm��򳇷bmp%�/����b2F��7����S�EY/��B�jg��'����L7Ĺ��_)dO��.ܪMn�f�߿��m$�Ssj�{�
[��K[���7Ӹ]�C�]�$�҅r�qf버!��=h��h.�|<Ә�/���F[���|��:���		$�����5�{��v߬69&�Ͳ(�s6��,��Jx�?Qg橞��H%΁��\��E#�y�Ԃ'�1E�0�3�Q��#S��g�_p��Rm����N/n�g?���r����+N�䚀��
�䙞(Q�ӹrq���||t+��}��8�lלx��u���5��� Z5���< ���� ��pS�����0�}(4蔖E;9�n_Kޅ��AT��C8`�#iF���:8&J��"!�ǆ��m����Q�FE_6�En�fͼb-�^��7�qA�?T���l�4����B=�����u�;B���]?�O�X)'F��$9!�f��\.|"h���4#����h��r2xA����(�[�}t��1<��&ݩ��0O�ƣݓ	J���l�ƉH�����pFewo"f�pRa���W��&_�C���B�-���>� �����I=��n��X�^6�{]s�DE���h&=Ŷ�����j���A�=0F��2h
Rs��e�zWze��6c��C�I�d��4*$kL;���c�{���s��1��r�I�#�K������0|�u'�.�m[��6��i]a2P�[w~ܽ����¡�S���1�݌K�g�>�_ N���[{���%F��j��(��(�x�"�������6�0��٥�Έ��_�G�L�	�fJ#������ f򪼭�C^�x4/��)�H�nd|cecs\�B�B�g����ǃ���˒X�d����s(t&b�=�o�I:l������~{שE.��%�B4ƫ�����N�焮�?%�H�n��s+�Rr�q
�?��|�s��6��Jd��ay�	����{��Q�e���LF�	�	I~>Yni(��?9h�珜2�HAX����l�t-�zc��HE��$��u
#�IѡD��[ ��f��5��&�B�0�;.�,��^�K�
�J>[�%Y	�t`�ف����Ju�&�Q�+���G�&�Y��U�t����Cx�9�t�1!۾����"8kW��8��%�y,H���O�����r3
��l1��Dkv~	��L-B��h, "�P_��ťK~@"2�) �+���C Dc�a踻�8����s4�a�����w��4�)���?^-�"�O��bd�f�{u����[_�Z���Y-Ow��G��!�|"M9#x�C��bBi�0x�^=T��T�z����TE̍����= �����4���Ԃn#�7أ�m�j3�����E)�c��j��qq��3� ��'o��[��g���.�w����.���^��Բ ��g�<KIʷ��~��� �ڲ�`aY��\�'jS0�Z��TqϹ���O%]���Y/y�J�$)�w��T���a�+E� i����^b�4�����z��~D��X�����4!5�r��(`��e*�]	^����u%S�Ț�p<Bʊ @:>t��X�/��l��?�2f�{��U��t?S�0Ǳ�OQ�{���"�%\՟;^��d4��A��^�r}��4�f��#1\�	�".^w��fv��V��@+�����R��2�#I���F�<��S߭������f���������-F��=|~�Iб���̤��ʈ��+$��"w[�^?.�k�|!��ʛ�흝�t���˽�� 5,gDn�sxz�ێo	�=軇�FU�_��ŕ��7NN���J �=�g*�̳&�ŏ�%�QA�}������'��o>	.r��65{?��fYh�d�tF0��?�lX ��ɶN�=!�LY���s�p��e=��e�ӏ���~�#oe�/�AV��(g�5�7Yfe�4`������r9��)�CS �*m}ZPgo����IM� �^:�z��k��DTlZH�yU�Ġ��i�~�^"x�^{M$�$�3��w'g6��?bQ�=^m���WḰ*ُXF����	�8����2b�@�#9�YĜ=��$��>:C���e�m�r@��k�>�-���E�)���#om�D�4��|Y�&�<�����Q�*�@+��.'$�)�O�/q���%�q��G��3�|rN2$���o�+�Ǉ� �ʇ�����2R�#���n�����(~Uv}W��@~C'����$��*T�O�-�uǰ� #D��+�U�h���z��4��*�>ig`�PU�ySH�~�~G!�m�C���Ӹ�P�n����һ�N)��g��%me�=`$
χ�p�C�� 	o����7��pM�>���+�r���z���0E������
IR�˾���!_��&�����5d���߬�$�rX��,B�i�{�L��G;8�X	QX6�n�'���T��#*��Bi�+��Y�S��;W����.��o��U�� ����؛�\��H�'�,j���ݖ x���ق#�jɱ�Me���]>�<��y+K�5�b4�D�K�y��؈��v�Y�;�M��}~H�PN�zN9�q�OW��Ն74�Z_H��&��\��)�˜;?;�/Lh@�� C�*\A?԰I�-�<�y� ՅW�� /?93�����(�0N�+�i�V�m2G^����b5�7��������>(P�]�A�t�^U��.F�=-��y[�O������+�!o$���q�b�8$�j�E�Á8��v��ᑁ��}�X��%�ܻxc}� [)MŁ�3J��M�C�<�!�����k9�~a��1F�u��O�-��p؁;��]����-w���
$%S,�WT��j�!�SQ�๦�<���D	A[	��\=�����1!��@���oh �r��t�!���RE��ִ��S�t_�D)���Y����2!4m GV�?}Pit��xi3��p�'����IA Egq-� �tߗ��ɜ���l��ŋLY7���e&JkӖY�p8�C��D��/�쎈�mN�B2ex'8]��i7s����g�mۙ-�"���uz��f�Dw&��ǩ�&�~ַ��,W�΢j��{M����Xj��J �|ɇ���Q|�!���T�?]�L�w�;/Nf���. ���Ez���("`���8��t�������jͦ�AJ�p��]�����ӷR� b]a)�YJ'�M�{}�%3?�������D��I�a��J�����>�Q=�HD]#���kVZ[9��:[�8��m;�ֱl��A��ji4��R���#��U�=��8�Bn˪/j;����%S����j�X�� 2�b�s[�-X�o��M�y~����0I��g�: Jvd{���r֨�C��Pz@��&����Z��| %]���iXd��?�NµUCk���=�EOm����7�����v�	�	Ђ�Do��}*a�hY�~��YhKIE���Ӵ�ٕ�P#u�)}�Pٜ�:��b��DMC\Y�hq�un�
� ��fW`�x��Ri�r���G���1s9;���]�;D�,"�l�D,�%�d�~��kM}��8u��~2�_�@�����'8���tf0��m^:M�>r#��TW�'DQtj�DJ�I�M�S�K�m�PR<H���hТ~I�CXu��[ �'������ۏ%��0#|�31��O2�p�F�
�����%6�+P�����O!V,1�ҒZR�#�����>�foX0q�rx����j��;��z4��i����@8�G�8�b�"(�����	����һ2�)�BB��{���G��aÿ��!�8��-P�ydTi��������)H�&�$�)^��O���
2qaX�0+'�Z�O&�U�vn��]�zX(?�C�H�F�rkT瑦���Y���폲{�+���"�C"Ԓq��.�l�l���a@���H�=E�ٓ�@��-pr5@0������?�d�����������9Xb�2�>�ݬ@�\�c���>� ��^}4T8�I+���'v��dg�DH�W��kUn�N������7b���j�����7�b�H�D @�r� ��rX��b����NUQ��ѡ�W8󩑼r�a��[�g�*[�$&�7�b�|{��"D�E�ua��E�c�eW�+T@>�0�(�wG��Ա��U��q`C�_���q�_�R9��S�ӑN�H0uo�*�n4H"�3���6KroUF����`��b�.�������[>�:!�i�ߧ+w�z���^Wu
e���14��x�b�v۪���QC$ǆ��xtA�W]�DTa�]����k|�q��M�A�@0�֝ɰC��3I#{�� �q��@I��z�v��V�����mM��ť�*�S�Z^��0�}Ҳ��ف�y�(,�p�6����������\����"�nsI���hQ�F`Q��-�;I&�D/����*��,�x�xɛ�����m%�&��h�G,2&�c��S�AT�uJ���=���]�K@��Q8q�k��]�v�f��mV���u�ވ��W\r6Y��I��s� �r����CM�����x�N�=9�Ň��[U�N[p����"��9VAJO�7�c����[�
�K�χ/؃!ݞ�(^��'5X{�i'�@H���y֕&h�+��j�:����8��2�[[۰.�0�8�	Њ����~]";ja���e��I
��p ����i����T���F�����.�t��i�Y!��\UКH3z;%����F#��$g\��)���i�yq0u��~
)��)��9a@�RdT�&�f)0���w��'��~o�dS�gߞ�t�K��pL�0�{W��D��ya�?�!y0:��Ť��y�6
���%�0���f7���Ƶ�L�a�,��v��V�a*�N�!���?�j�k{tO}�۫��oq��z��G��U���"�j����,?J6�s��V)D���J�+,,g�4�&p�q��=(��B�]��:$�h�*��ͅ	O�̉b���+���^� �a�!��H:��B���i�3�V��)�c���l��\�3[�=�"� �5baG'r�x�Y���Vt�T�P
�u�D�,��ˁj�
i,-�TQ�0������ty}���2Px�gl��7 sa�Hn<5*����D�Ҧ�;>?��G�e��J�����/����w*k0�Jk����@�J�Ф�r����W�u>>ް�p�gǚ�;O������η��  ~Lr���l��;�-*#H��7s�F1ǖvI��Ϯ}/��
�����˗�԰}L�P���W�ak	����*�~M"�ʴ�5�T�Q�X�8`��"�jN�������P9=���se��Ro8��G����,4����]������l�v!���:�;���	�7�m=z���*����|n���2�����*6��և����хשI�~%���"��� �81��+��e��$��%#:���%i����s�U�
�zY�b%�1Ѧg�-*$�@�y%%(D�uu�0�����|�#��r=���eJ8Dz=k��@�l��AxE0<��EE��zz��6�)�4�|t\1~B���2��_���+|uӺ��3f��xx5
��s,�Ժ��l��$�Q�x���o�����~c|p�<;~g� O^'ǚb�l���ǯ����f���{��;7�{�A�:D{Q��x�#��2�T%�%R�vZ^�r���Eҙ9����`�B��`��3�4`:�e���8�7�|�<f��	��?B䠮3��;B����2dE|�0��$bQ����\�B����	�l�q8̬M�~l�T��@Z��!�r�ΐ���]w�o�����;��<�����3ԩp
�¥�hx��tM�Sw����|���:�K;s<P�r��-�$nd�֬fYRg�%������CS�������P �Q��`o���@V����T���#Sh���T��K����3����;-�vR銨v�݂Ù����&���������0;w4��C�n��� E��ahxD�#Y২5�Q0�.������"����j�D���=lT�L ���K�/$ߢ�=q��wu�0�N!h��r�
��_��W�	�7þPY�q�b/@Y�\�H-8���5ļ�tj���<N�i������� �#����(N$Ë;^'D
��+����Ń3\!;m�C%�>�W5�-=b!�ޔ-ܽD��1q��4�A[��}:��܅:n2�0v��6��u�E<�A_��f��U�RL�F��^��e�X��3V3����<y�q���v ?L�@T��-($an�:'�mʯc�B �V��&��ev�tRv���)�9(��ҮUR�ܷ}/2^�]k^t�E(��L�?��mv����PH c�A��0�$�W��� 
���Wj�9��C��M�VOW��X��X5,�*�)�L���4Z�~(?Ş��K;�����n �[�X����,�47��D~��:J�da[X@�kU�坥�
����|>f/� ��3�r�;s�c^D�>��	���t��k�tS�ƅ�S�6��J�4����� ��̎��Ҧ�=B�혂�"0�R�VG�r`�(�����F�V��9[l ��--�[,V�ꅠ2����,{��Y�7� �殺�ש�D���q�4�[f�"]6ד�+�GS33�*���y@�
�޾8Sf��$��k��)�I�m4#n�1�E�Ƹ
0prBZ+z��5�Y2��a��į�cl0^1?���?��ZJX*}ְӎa�2���֞�Q��/�f���{��R��?�����s�y�?�܌�����o���ɸ��'���JJt;p_�c3�HD	��Zg��%lX�2\�E$�y���$��P�T�'_�E���x�+�<"��1����ת/B
��ZB��� �_�J"6��q��Ɩ�� �V �������|�B������ӂ_?��3M��؁!u:р2t2GԊ��Z���!/������-�P�0Y�څ�Ax�7� �<l�Cǔ�h���H��iZ.��#2��!��Φa|C�߉��}8�_0��9��JK������\����e�;�Wv�M��^k�쎈HV�O�)��9�%�{�l�b������}��r~/��G8�jS&E!n���T�޲|�n*��x��ÀU���`w�;�,�G�m��@�"D{�A�~��?�;t�v/�g��V�x���l��EQ;O����L�l��TM� ������I��$R3��G>	�w,�^`�ӽ�;�}CL2��8�s=�#�2�ʩ�"��b��,k$:��Z $��l#:V����IاI=����/s�X۟�� Ү��,]A�0�ΐ3d�IV��;�6��0+"�J(<&�8�����L|iO���X B��;��y�IT?Z%��� ����oόq�?�q��ч[Ń_��3���pP��O�� 8���~�mW������l��6R�w|@/u����i�:�h�"��B��b��vH�&�s"ŨZ]���0HO�TV��t;�I���G����PN�1�nS!���Z�E��ǈ�&�F�BT��۳���dP����l-��>�� �s90�z���L?^Ţ
�L�А�͊�X��s��#���;/\ZQ�9���(�Nֺ�K�=2|��Mй��V�5xG�S��� �w�Fq�T�h�߁;U1!i� ��� 7����.ؙ�!�|�bԑ%5>`8�+���;n�W7��	������Թ�mU���ڂh^@�;	����G����9	9���Ƀ��P��]�����G/T�(���6닸��$�v���\���0~de<Rt�]Xtp%����hZ��ʆU����|;��i )v��xၝ4���M�iqJTv�^�\*.A��lrz�u��4�E�I�@��Le����d��%7SX���{�U��Zs�,�����T�G��䨯�v�ۨ��| ��2b2@敟�l�aI�Zp��TmEN�~T���{���&w��ч�|�j+I��;��U�8���woq)LW�q�����޸�0�@���Pܖ1���a~��1���	�Ƈ+׵7Ni\$\1����/��G���G2�WD�Д,��9�Qv��Ss@���V�*�Nh�U�z�ع�V��{NҖ�Ȏ|,Ӟ|�*DW�臊��2��wW�L	�� ��̠��;OL=+�� �VJD�B81w�M-]�z����Cֶ|{�"�,J�u�I3����<��U�W(�q��|U�(��9� 	�T���}<O���T�Ȭ���fPѢ܄:���>���!H�G������s�c	���4	��KYX��Ü��$1�)��4��+0��&���"���HL&b�<�����GX^e�-R-��Z�E,Otc��<����E!�M��T�&�n� ���rP<ٞ��񵙘M���	w�^�=��͗�+�#
�r3�s��'5Nc!���X��z3��uݐ�S"���*�rr����~O+�F^��A�@��}&rN!M/��ϿWZ(?�ݽ��^rD��.�F��«�A�b�BgTYG#_V�<�Rp�#E�K����}R�%�t�	|�U�$GL(�"��꜎�v�{8�nd�!6�Ù��_�&��5����ؤ+��L�z��8.��]���B��CC )-6�����g�ͫ��*>��]�)�I���8��+u�$��m5F�@y�e�g9te�CU���Jo����щ�JΗM�<qc5����nkq�R������I�Z�(�6��ӧ/ߙ�a)c�6�Ś$K�UM_?�}�9~G����U�z�h׷u�j<��*e7�!��[O�ͪ��/մ~�mr*�aq1pb���]7] �X��l�)j!���|B�N����1��	'ɽr��Z[5�x�J�F.5M�x��Dj����jwK4�T��9&�K��x�#&��I(sJQ+���9�s���1z�* b�������L� ���3���!��A���|��[�cD��=;e��V�xpOhnX�m��@�Q�ǽ|�t��MJ���J�z��1�ĸO�wӬ�n�>[srCt���?�8j�D�b�z�7�B��삽��mɺ�����#�vO���Vק`���<t���j>-��mw�B`Q��`�:�Q�;k��d�g� �m�1K�w�0N��j��)L}��8%
~�O�kc��D�z1�x<��a�t2�����qKp�����; q�gx�A����@D��p+�ME���o�i;U]�
��GT5��f�݅9��}�W2��1�E0o҈rb
{KM��[��;��V&5<)/Z���m��Ja@�Bm�����ez��èڸa8fa}~�'j�1������k��޻?^q����ŭ���)��ewm�+�!J�z�o�η��	b�7�@W��FB�K|��6}�N�6:?�� �A� 0ru�Q)�\{�EY�v!��a��[R�]�(�v��2��c5��,sX��01�3��`�Z=������+�
:�Ib�Š��u�]���j{)oE�m�:��Q�\&B>d����t����5W��;
{� /�@5!K�m�d>�`�+�2�ʼ�jl�]�M.�}��eK���,��mPK�.#�ry�lw�FP�R#P�����\pF�Mt`j���qO��w9�%��b��2[Q��R��(��T��D�=ʳ3,�K�J�l��7
.�1xB�LC��r����:��~��=�-C�0tj�YiDحC�wM��g���A!$"�0wNh�1���F����a�ǈK20�~�[hܟޞYk�X�F�롁���:)���n)����� `��D2w-�����7$�#���/�Q @~2�w�Ҋx<�a	ۛ�Bߗ9b_�4{lb��B �SAd���!}>z�O�*3	�@7��,$�	��cj�_��{8'���;��Z�q����砠z2��Y Oy�/h�(���~|�3��+P�ۧ0��$`��~��Պs@���˯g
U[S�-���&����R�F�{Vb�l��4���,�mP�ҎdCW8v7�ݖ�x��n����~���]�e;��r�����[���	T�k���kȊ���fm�U���x�����
��s�@K-���@�V���Ŵ��my�uCr�XZ��ACM*W�gNx9ej�Mt�/2��5�uW_�TKhM 8H_�ج~Ԧ�GN�}r�|V�H/�;ĩ�)5?�I�V�"�M�ɗ�5kahޜg�w)���n!Y���E��}-�\gdS���¼�ҟ�_m*Ӂ���X���Ga\�P��j�%yF���i��{#^���${�	�'�n�1�8��cmD�(�9Q���#6<�Cx:��w O��lN�U���o����=65Yoj\
c����(3j(Z�PGr�:���K�qfvsp�ps�l`Or���9���@�[��V��<�pa�1C��-�~����0[�f!"+~1u��)��E"����Z�������$�V�#KT!��ͷ,4��+(������I)�~�M�"��mg�Ʉd3�4�sT�1Ʌ��^H����̘�^<�׮��97��?8Ȏ�,���!���������K��C�w�4;��^Ƨע=��L�~�E�b?jf3Lde���(�KgZ0'|�ė���Z��Ʋ��t���]�&Vh >4�㇁o!�D���°6��=� ���1�W;C*���YK4�!:����6}aG�����m��1�ϧUY5$�����:T��VS�������@�Q)3��V����>]��	�Bi{�n�9RV@_��*E#�>�T���c�U��!�L��~X)��ƮZKC�|��&�<I�,�Z QTэν#P�'t�����\��1yz�9}��jb�6���`��� �ʳ�{��g)DL�/5�1e�ۣN���ӟ+6px�H�6�~u$,�2��A� �)���dr��o�Ox��V��>K�� ���G??f7�r���R������X�T���<Ho'��c��EpKvϙߥ�Lo��9�����υ�B�J��Ula.�Ū�ڀX4�F�3�J���G�W���P�%�R��_^�x���h!����GI"�[^���F
�羢p��Y�I\�[���J�f�j-��x�v�=��S9J�)������7Ek�����������C�7��'=1����U���E��`d�UZs<�7���r��,@���k��J��9���2h�T��ֲ}��� #}W�z��%���@�Vwe�{o5�t�WS�T��7�a>S1�@˴�����X{n�t�ЮTmg{ES��.[U�(�ٷ���d���*�3��+�lFG&L�u1�%)>7�ﴡ�=�	vX>�/B�����*�Y���C��Zd��y�ʍW�ǝ-� R�[D��k��^���N�un��:t��>rfj�l�y��p{�{k��~��2��q8����=6M �G�:��T?�ᾗ�ǧ�L�G��/��h�;�K#��B�U-����[���o���\F��]�}ؙΜ\dh���UhHt'��d�����C��-�h�~�\�ե>����i����U���v��v��7$Xe~rGO%�>�D��Z�hq��pg�P5���v٫�Ւ'{�U@|}u�LC�����+�u�����qk@|���tL@��کE)ю�%1Lm�v��n�9�0h��TC�1&�H�ư��!�#���.x���呓!_�� \5�T���X{��	ց�24գr�������#u�/r�4��U^#�eId&�sY��*V�<k�l���TJ��kV��qjõ{/�Uؘ�ddL:k��72q�ǵ4�{{�F���mR���� t��乕u� ��]� fn�.�Ό�$r����<,oV9}8>�[�K���}��ᡯj����"(/�r��t$������a���U�������@�d���3Co�e�eE���p�O�2S۞���,�0�T9�bJ(E]�J��hh�b��\O\�/�Ղ�L����L���B{p�Z�(o��P_o��@�������!";ɗ���@�͞�g�᾽��3c>jy4�\��O��]K���t3i0�^y��>����$�"��M�JQԉc M(�_~��tۉk�G4�[�nz+XQ��t?[�p&�M�.�[�l����\I:�U�n]	&\y��4�)&|�����J0Ot�=h�-���ll��9�4S�����0�Æ�:���+��ބ;��@��-X9�
])���,}�;��$~�?�~ʐ7���J��L3�g����x*�U'l\H`La�8aL3�/�ud����l�^a���Y�ʍ�*E�;�Z_ ���#�c�������RLV�/�0`�?�-Oϔ�J*<%P+��wX���}w�ⓣ��>�CE�v� dډ�/�Y:�l�=z1������(�*v-y�i�#�;ԣ*ϕ�_��d0�'�42ۏ��?��|�̡~�����B������Gri���̂�J��q�BC�T@��F�� E&���\�|������+:�P+O?�	Z���|,�ׄ6��<ʇ�����pw��@Of�y=�ȿ��Y�Hl�|b���8���$����)�[ps�%Q���)��D�:��?H�3MzS����@�V�`�}���K�*���%��_N����!�#�KHu�'�9���ٮ��q<K d�h�0t��ar�(����;`� r��R�fMc�?��B3
�v��n��8@i"�n?��j��)J�@�G5�|Ȁ;����m�pf (Z���fH*��j���ݔ��+�1>�5^GDXB4�����-~��S���ܫ`�$DI׏�	�F=�H@$HjH����"/�
܏��>$�+�-�=�2�aP��Kf;�t��P��J�İ�> ]g�C�
�{��bI�)ܯ���r`Nㅲ3�3�g	5ڈ�@^=�m\pة����J�u�Z�5�G-��� �5Qc����04�N�5��\���S����K�U��L� �gZAn9"'�/ +�OC�:���h��ͿY9-�N
?9/���7@#@ �����a2�&�@���ŐƗ�ƫo��;�q�j�<���B�3��V����WT�6��ҍL��+�A�OȲ��u��9��p��t�ۊt�����+��mo�vD\�2� �{����B {�s�M��t;��Y��A���+�3G��}���+t��޴?�fps��,�&�����&%2�Ҵ��{�@����R��wx��%���%�Ph���Gdtq��(�1��Ap����~X��	�� �̣�D��a6f����j�3��m�[&�1��<.�r6�RiÃ���g�țq<Z�}�����b(o���
�e��J��G��#��ʽ�ʼ1��}��TBߋ#|:!�y��c=k�l�@�7����RMFgZ��C��bT��r:�G��{����y	�,�wQ/Яކg�j�)��eO(>i>d�$���̙e��U�/fYOh��.A�Wȡ�&�1Ӥ��؞xmF���&?3_��" 5ҹYgt�=F��U���dlI�K������
D����q~�]e�mpF�w�V�����f$��}���쮝b�ѱz��S�ZZ�ޯj�~QY�7E�F{���[0���Y�����}��u���� l��~���+�U��Ux��7kPWk����lM�b���%Be�x��=n��p��� D`�~�'ކk]�e>t�	�+Ɉg�E�1-��]V�zgW�� 5n%e�.�埬rs~�B�ySs�w�1L_����8��}c�q��X��B�[)�u�D�<�|-��M|�&�����8w�q��)
���Dp����S����?9�/������y"d�h�g�}��; !�פ̇JS��[p4R��x��#.��s.t��o��u�m����vd�7��m"v�5e��_��,�1gw�H9�#�������_vծ%B�D�Jx&Ӌ's�B�=�J�L�����vɨx׉���Cw�tA����p��{��A�9U�zdX�To��Ǵnt8�I���9B��	x5C�jG�"�k[�E#-�!�o`���Hǂ�)���!5J7��;��-�E��_�����ѡ�����=U����1Ɠ�!^u��_鉑��3ܨ�p�V�	� vK~�j�����u���<Z�[�=���ā���HC���/#2=wr��㛯��Q�1vU!
 
��ݚ*[��+��]I��C�vkRCS�� ��^O��m,ū܊�9Yw+�'@���߇"��6����f�zd��)V]B܌o�T�ȱ�͛E���t�t`B湔j�J��>Y�:���(6]�Y��R>Mj+���q:-��W��!��tyj�AA��T�~>�2j�\b�T�&a:�d��7q��a�r�sf!��3�V��_����� h��A�"{��s�
v�,Ʊ*�J]<SJ�b���!�􏎕�)(����9�7֞R�(��xқ8�J�rA,`���\��+���(U0�W_K�2 �J&}�"�������avw�!
�-�DV���ڸ/vA�\�B㐇�\�+��ġ�
D�����g^���o)�3���t��u�
�o�$���eG��yI)�H��=M�Q,7���5'p0�����fj����@y�PMk{#O�+A+�����R�}Iu^ҢZMo�b� ��#��םHS�g���:�A��>3�30X�����@�����l�ha����b�i$Z�bB���3�F�{�D[Ry��k��t_M�ʅ��f�s�tVP�i"x��w>��o��pj:������+����������
�q��������B1�o�D������\��J�w���h��9�r}!�V�߽_Q�I���7��2���6�p�H�x�D� R+4^9����$�<���
���6n&�KM���u�G+Z֎������Wג=�~%�;�i�|Z{�w>ץ��i��(�X)8M)��ǃ^��H�Z|Y_��}���}��(]�������1&�a�p�%���F~�j����b�$X�0�<`)�vy��D�E��"G*��T�iq�^L������ë�DF�@�4q����{̓=������q���N٪lY�Q<�W�:k��Om���s\L�)���v�}��^u�:r�:c�H���Q�\�&θIE�M�H��%b=he�O'	�z�Ѝ�^�����KMk�X/Z�S�I$��X':|��ڛ�_Ci��@��q�t|`A1��
��9�~�	����4�Qo�r�2?C{��Pp��f3|�L($諵�ڞ)ZL����-]��z���dR=a��Z��+kM�C�y*@��߬U\+�&���4���n7���o^u�&�'�xʝ����P�N~���U9nή�]�� ,�#S�\����T�%�h�W�ëU�0�|�ߑ��_��"F6��k��)=�$V��!�~k1Y�jy��e��������/��@��b��~3<7_ϣe]n�	j�2��c �Ir0@���%ߑ���U��i���}Ix۳��@\�ww���5(��kU����I3��vZ�ȧ�?g(���٧*58�Q�T����6�n,��p3O�o��9�<��	���P�2R�Mz��N�D�![��G� �8x��������H����z ��)�Cb{���{�ӕ���WTX��*��ђ�pݠ��_��E�h��}մ'�ñ5'���&@c���#"*��
r�?�.�t�w?A7E�;���}8H��By#�{��o5�#༯!nn��;�^�r����e��Hȭٕ�^��F�H���^4 ��J�1d?E�us0�<�;8fG5�ZU%�������8-�gn�|�.�f����4D7bB�ԀJ�����U�w6�2HW>�X�aX�2a�t+Ԥ�7���M�ڋ���<�P+*��LN��@dɳ��-��(�e֮��c���f*��d�qQ�x��X��p�Q��x�?f7�Q�n��'����o�Sf�ؓ��I�D'"U�wÈs .a��>^e�M�!>
�2 [���M�^!+���ʃ�������D��}��Zg�Mހ�,d@�Q����4�U�3iV��^x[϶��@ O�$�LؘX��G�*�2힝x��L���)W[�֨g,Ͳi����t�i�	sS�~�"��ȓS����X\��nL���Ķu�K���
;�2�ԧ3�/q�]\E�s�q�'���-�?��X`ֵX�{�8�(?e���>�x��9U����%q���sL��k��n��u�-+[2��-�������[���>�Z̮rj$\��ᛢX9�.���>��P�n�YNe
��\���~�ɧ1��]}��A�Z�H4��_��?(�~�m�j��I菾vҰ�D������CZŕ@�^��O#R�W^ژ_��aY��N�Rd�?��k�
F\3y�V�����X=!=r<dT�Fy��(�7:K�ȧ]�����������l������XǍ���:_��[�3�D��W	�@J�����,&i֠7�y\N�Z�,>��B�&�:w�?$�_ŵܘz~�r0����I���w�#��&��.�um��u���s�j���Y�zS���g��!�Z�1��;1q��96��;�mk��D�/��ظX����ĥpӠ,O�D�.�.~$�K#�,`�v�;\'#�H�F1`E���m"��oT	#��:�9!��q����iF=g����6;LY?�XI(C������VС�_A���K��%H�~R��.)#v������<��.���2����넷���Ъ���xc���O��ﺈ�Jj�5i_� э-o"_�����(��*��ֈ���a6�ErQ��i�~yX�
�����~�c� "�h{^$� �
�[���F��n��Ƣ�<f4��I�zX�ӏe�iw��wr�p�{:���[�o�O��X���E�^Ss�� SH<�JuŚg�S�t}⿶�p%���JrL�M䋧�GNV�W�-�)�B��қ�l�'�%݄��;�"S��>P�heg$�Ĉ�=��&q9���3^L���L3o����6��`�"��:!��XJ=��Cz�L���W����GG9�ʘ�<�@�R@���iZ���$��-A�tRՔ
F9��p���<��+��%퓮˔3��;�z+ %9>��Q�d����� ����@�㘁|Q +��z��XHڣ|���z�m�������lIOK%���}�b�������1�mj9�/<%Yp�"v�H�'S:�c����z ��7���n+[�|��X�}��,+�@_�_¾g liNy�B:������T
�j�?�B���O��+W���"s��7�1����@vFq��jx"��잔	�S��|�A�s�Hk%OV�����|��ܯ�j��-��4l�H�9�JL5#Nx��k󎦚 �gݡ��¤�)_B���Z����W��� <��Ŧٛ]��.	Ng0_ܵ�U�2���S�OkL���0���;�d�a�U��d�o ����\̙9I~�6�}P��"�G|�T��LEm��Ug�?�AJ���e��ye���\ǞF^��:�
�	�ki(�M(������=���k���w!X���U�c}��ȷ���rR�;�E�-�pR6l�l4:��50�T�bJ��=���J��:1�A��UYRB���C����+�ʘ��V�����8H��b �ʴ�����b��J[x��sәVm�*�P7�0d.�bd�F���Z�:^��f�\��U][�K�Dd���ә~�v!����	�6��|Xnоh�V��$t�"���悁nR�%V8$Y�t�l�q�>V�KUP���1Ă��� ����#y��-��̊���Ec��GQ�B�Is���!8�x�� ��Q��8!���b��*w�	��a�����TȊϚ7�:� 0��D��y�ͪo�Qw��kO�/4�KNS���F����	�z���`���ڨ��,OT)o|���#р�W�'�4~h�K-�(G�Q/KHqe�5��D	d������w�f!2�UZ;MR�[�4�)J�[9{E|W��c��n���30+�������*wC��r�������Ӎ�p������[�4	��B泷Im�c^��)�V���jQ}�Щ9�d�5s�P��6+���l�J���%����fM�.�>����.�a������=aq�5)�h�X���jQ��X�4�'��_ڛ[s[1Ҡ#H;z('R�۩�M���v�[�m.X]>�*ȴ6r�Zɒ�H���ci�@�����ʢ�(Є�����_UB�jT��:[+��g�4�3|;t�b���eAW&�Ա����b���pj�G»�� �#|�l)qh�ʬ�^�I\��^�#�?[�_H���P���4�p����Nj��򘸃d�V7��5^�tkK;ެB/E��\�ʣm?��	�j������!��4����x!Zz��`��q:��ݚ����W1���c��Ib[�T1gא%���'§?ؿ~�p^�E8%�Rsh.���b�Co��7Z�Gڗʮ��\1��(%���~� �±W-������@��y�@f�e˴�~AUU���V�����g�n�RRh�YA V�~��hqY1^,D�}�6c,�M���&��S��v.U�cu��8dO�s:�c� u#���
9[ͺ/Nz�����ʺw��Ю��#�rqoz��E��w��F<dD)�{㛧��:́�V2�h��*�A "�r#��? ��f�<����|@Jy�� /_��akN����}pJ׮�с��>A���M(�������U�FFB�`"@��S�K�H����B`iI���v�-��m����P���_�}���1�ng��XL�S��Ń�Tw��\�1�1˙�)��yE�tj��1��`��k@�t��1o^��з[1k(��!u�T;l��C3�Ԡ*[�\iZK2~Y��Σ���S�\�Z�E��gd �e�O�C�D$�
l�P�mO8�5��N[�ŲD�����j�h/Gz_��`H�
�c�����a+p�|�N��X(sSZP�\F,A��h`�1�Dw�k!.�	��~S=-U"Q@P�C4�z^y����'<	�"��q�S��\\���T]l�Rg���=�{1lh�����n��'m��v���u7��-�H6�'�_v��>�f�[Z_S1Y�aP@�\zA
G��_��("'B�#���8:�'{m�ᔷ,5,�"�^����_�pm~�1����ުF�ـ";f0dI���^����d��O���u⫭�v��S�Kz�.z4��p�.�K�h�b:�6@LE/�ȼ<��à��7��ߗ*"����X3ffc��إ��]�a�n�ROc�=X(�`�	����0�"*�)b�A�R�˶P7�-�|GB^�r?�l��Dd\����r?��ɯ�Gj�d�mudYX`�"�Rl!ì�������\����{q�nl����Z#:�ժ�`�U�0@2������P�݇m��l<�$s����P����0�F��:�k��� )�9%�6�d(��ɓ�Nw����[�VBԲ�*/�WtY��W�?��e�4<;��U��-#��XRl&�����`�>�?��O�ˁ�ݙ�'O�u'���G��T�D3��މ\�~`ToŚ��ؕyF1�}2T�D�>��.��6��6�X���D7�dפf����Y�\Q�,r H4=���(��uy�s&���=�{�,�gE�8q�������~�S˃�5{�'�8/Z�ՙ4iRG��j޴j�Ɯ����4Ɋ󼱵^iڻ�>��oZaɒ���`
�c��`�k��賴�Im�r��e3�4aXQ}/9t�j7��S޻��sS�j�/ݟt��|y����f`�2�!�Q/_�<��\���&D�'�#Hb<��&������;�F�VXg�����g�"Z	�瑣�Z����{�)��;�P>1f$@�[ŕ���]%��4	���[;�~��z����Z H�X�3�0٬�o]�[Òj�ZCh���N����a�2ihܯ�bzJY���M>Ɣt�N��I�a��F�_�I��s�O~@ې�*�+���{�c�S���b�@��[3ݡ<�jk�n�x���'�=Х7+�n����}��Q>�"�\�\Š���z�<`~���![q�����%k&G��|-V����!���W$
�q�L��x�!�՟ft���f��_'m:z�M�F�R��O���_�4��Y{2i�i��/gm+�?B��F�V@���<@n%�9�"I�k^��jk�N>�y�%~3!Oo|����%n��i�M3	$�4�,��|�\ⵃ�윅>�f)�uĜ���Fu�?��T֬�a7$��C"eR��	�J����@�������=tJ�Χ�3��я@(�{H�`��}Rg �&���M��[Π)ȯ�M.�T�	��|���%BJ6YE��PJ��5#{3���i_�4�l6�40Y���̫rƇ�� �_����#�#<;�~�T(�s�)� �BCxy+$��u+��c�zX���B�Pu�}�F<�gvޛ�Z��_�~�����Z%hg}M����6Y�J0;��H]��?�j��f��e7�Y��'h�����P_w�<�C�F�3G�U�{ �H��t�>V����J�����>����:Qk�\0
^l�5�}��ٟ�Sh�2�eG�З%�,7?�%y٠�\�q�5V�p�sp�|I��D?Y=�*>���κ�M[�� �#�I?(���u,@ԯN����'��U�mL2�7��n��s���O����I�z\G/.g ��.}�*�Yi�+5�o�.�hxE�F!�{�?bE��[����)����T.IMpw�W*k�g�pM��i����8������01p�vokh��x$.{aBm�_X^rNv�'i�s��⑲�<����y\�Q�_��߷F���>��yEC�=���M��� &^<9��W5�#벾ɘ}6��b��tT5�)O,�������<�L�Z�T�C�3�ʞ�֧�6c9����Y�u����ʄT7�-	�eë�&E&*�U��j�U��4NhdD)k[���|�kA#ϼ[��/p�ܯ 
�>U��`��r*�d�?L����s�m �*�*�#��	�D���.���ݲQ��soTT��R�97�ᯛ��B$����f�y׀x�쇿s��2@qm��e�[����#�R��7���P�$���Վ\(��Mi�����'��g�=K%�A�����vHG%
�9��ɿ;��|�u�7�(}QR,������㽪/#t�nu�ΦJW��Q,�w���U`��khT{*c��ݬ�Dk\{YadW��)HO(yq"<� ��?�JtU��pY���l��Ǎ�D�R���� �*E�RD�
~�y�C�ͳ���: A�,��T���V�|S�2wI8�MvkF3��0�GW>y�9��_�L�������Q�I�G���5E��˲�K�yY����46�$���rk��D�aE����~?�%p�j���}���B�%��w�J�W�������8���+Z|_b��X�$c��'���� ��
��j�,��o��;mP�����`�ǫ���8˿DP�M�ʜAG�,Ze�Y�Z4�g��5,d��IBB�k����GF����/��
�)���⿹�D&s�k�ҍ�)���2|7��q�c9�7G�����qJ���)�<��wz��=UBu�),g|�Ӷ�N��=.`��i�Өa� �w����4/�sI��˚�����O&��O�/��!2�#�Ը������@�I��Ĳ���nl%����ӄ�� F�ej"Ɔ����6���K<jS��(~*Nre�d�<
�W�Ig���O�a�G?�vE��~,�k��J~�� �`S%�3�I�G*a��%��k�m���<��m^�g##�)G�nѮR-�lf������R$�F�+oH�F� ��.����y�
@��Q���%(�w���[K1�6P׆�},fʸw��zeMH	��y���S5�#��a�j�Օ!�^"љ�ta�=�漦���~��U��gJ�?I��Fw��Lx�D�G�v�řI2��|�&'�G5��u����ؙ�d_c�@9��w��)M�1��۳�z1-���3��{ �˪U�󄓠�"�K抖Sh+f]kq���?2giƴ�k���_L���w�/��y����^��F����@�z��g�w���bdx�l����8�{���.�9R��J�ʡ����ݛHaH�r,IOTzN$ß�3B&���&x�Yz��Y���\�A�,Ѕ���n��%���șU^��~,�&Ӯ�q!�Y���Y^�"m���x�V����3*��|�O�'�u���MƖer���8�Oe��CwBgeE[��iJ���q9�v���=Y����.=M Q[�ąe������G�+xVI�_!��VGu,'����Y�Iu!�*_��Y+B��BOLZ�[�l�$7	q��2g/��(��aFq���G_��Ք~x&u�p�KW�ZNk��p�����qM!9�uL��E�[wqB��a���52�.�Pu���׬�͂hh���Tw���Sn{֍�X��N=�ˊ��FS��TNlfڿ�J�0G���E�*�*߲޺����J�_��=��wN7D� I"4��Nrj�?և)}�*k{{h�ׄ�|�6����˒G��ϼG;H�Pz���:�s5l���'�h�n����a]�T��fLv�eY�SSo0.������2���;�X��M����hb�h���wIz�L���C���@���ӳ��42�e]���==�����9_ύ�|�`7�E\��)cr �L��1o�v-�zZsOF��]��v�ye��F~2{;?�6�!�ݘg�IV�������c��J�\eĝ�gC
g��I[K�=����"���, ���m���6m5R�#�6�C�+�8�� ��}�؀�٭/�O*��>�`U��Mu��n��X~�o�N�m�և]� ߅o6w0�9�_j��n��Dc׸�]'Ү�M��T�5`��
4Ϝ��ǰ�;���b�����U��S�A�Q1�l2�cR��D��&�Fi�o�F�W��@���\J��eQ.��JS=�*"����@S�l���� 	uU��@F<8o@^�\��)�8}tyU�%	5܉.� �εcW4�v�>�~ƌ��}k�l{�'"��]����OgXg�DӀl~`1w+r��D��������,�(e+��s�7x.�V����Z-\�+]��2�~+P�2�j��.�O�1��۵�xٞ���gr���X�5*Z�����f�Y�N@�6�l-"a��)rLK-)h�����"�rV�]�[�$��"S�Ce�.�
s,�9�����k�)�k���.$��^�����Ij�Q����?l�!=��l�;��D�S��D�Lv�A�t�fh�\�_��J���S��p~������5�[Y��ƹ��}F�h�-m�|E��^-.�o�R}�)���~�2��F�HD��bQ�Ʊ�m�d��j��!5J��mL"1}p�혞\��5O-�+�W-"�z��BR����̈́3�W�u$��-Y��������Z�������7�
t�&��kP�K&5|��5LEG�k�(��1�<��V��T���
D/���P�Ø+p0�-�[M�OYNg+9G�"Cz�j��Ө�dk�'e�Y�T�W�/� ���aSb��v�vT��V�����mUS=�u��聖]''"����a����ի�L�Mz�hASFU�4��^��y������ÄP��!}ü͐
�g�oe�y��yY0 ��q4�$V�`g�ǈ�~��2�"�[�9�N���|y*xH��@�䜽T�%�(�Рn�&}�}MS�Z�Y�I�0�O�蕟���q�X��s�EBΐ���u�h���Ac%�3�v/����N����T�U��"
P�ɷ>K~����?3�E�:����Hb�IŜ? ���{�GʞU�w�G�ֺ�s#��oo(�����d8Cw(7c����eK������X��؆�k�g��թ�]�Re�+�$e�w0nJ�"k�e�R;���2:�;hS��i�`����j�����Y��=h/��5H9b�D>ڎ�נ����VB�Gau(z�F���yZ���+�]˙��^��d0�|l{;��87p��r�}?�#�����zN�`C7gX�O��q���X��<(��S��?RIR�������2��#@�Nz/oֽmQ��YhGb`J&u��3�Hwh�+H���u�&y�?�o��Zg6�O���A��A�����Ca��<��UFe�v�x�=E�R�oI�|.�C��[D�l�US��o5�!X���Z�.�qd~���b�Z���mO�/�wa���gRfBh��_fGc�Z��JF�A���S$��žz�'�v��%؍en�'/�kpT�<�ݵ�jY�D�-��z���p���7���L[O1�mx�<���K�iÛ�NT9D���u��J�3�$�]���V% �KJ8����n�������dbO ����>�N��3��LJ8�A��`P�.�Wj��-l=�mHS��6��G �w�8;aHp�c��M$)����*p8��K�{lzoOz7D���i�<@�O,��O���, �T��<�M'��+C���b�E��~��߽�8-BA�K0�$�j��Z�Ό���\	�gV�U�]�j4���g(+�'���*��"?��Ro��K��.�|�7V*�Y���߉�j}%��F9��JiǸ+��T�����A����
\L�w��{���7n��ᒯ�y�)&�_�o'�(��T��M�z�r7����Vu{�~o����"�lŒbD�[����`G�j�� �ǁ������"@�J)�q7�bo�B����; ��p�*
6���I���2�����t`��!=X�r���k�-����x�ج�km��`�c�i��+ɓ�?��z��2�h�c���P��i�m�#������ZL��6�^�|�X�űk^������A����`w�;�o.�}��4��W��Ѝ�v��v��=����|���T[�9i����c���1�f�6iDޟ�A�&�2G��1ؾ�=:��U�x�s�SZ��)g�%.���n^�(Ĥ� �:�Gɘ�@�Z�Ϩ�T�n����Iv����B�B�y`D@<�����j�h�3��|.��9�m��8ݼ�c�c0�q�[�0W��>1ɾ�+::�c����^&ٮ��BV�Z��k�6?V�/'�VK������I�6����c�$5>NJ����2�Js�镜`�1�d��u�}�A�����d	�"���Yf��q��K�69x�,K�g�����K�_W����҈ ���V�����yL�B�ބ��bc��'�Njc�m��@E�G?�I��쩉c��eT�6	#�~�e 5ŉ�U��e~����2�q`�zWUZ�#���^X��=1�k�ȱo	�����c ����*"� v�G��cO@��96%zP��S+�\�ޭ�ໆ��8�,�Qc��|:n����q�~׍6��jrE ���jChܺ٭�3��?ѩ1|�#n1 �Z��Z�YI�K�4�4��o&����ǋt�qjf_��04���H<f�}����ڇO���2�c�ǡl����A��;l�������A�}���
�s��D��@c��!Ip
_�\4.~E��k9��`�W+;�^�!�F@�=!�a<+��Ŧ�z��[� R����� �)O^�z]R>K�	��#߶}:�����<��1�R�����>��11����4f��h��b�Y9G�fl�:2�hw~p�!!����7d�����Eu�y;�����[�/D��h���^�d�����A��&t=2)��{_h\Z4��-l�;�mG𿴢-$�^�2������D�$JD��
�->�i�&3�sӧ��4�@�3�-ڭ��ǀ�9!�mr�D�c(8��0[CߺAX�F�F���$��e[9���_?y�Z| �>��z����gFr[*Ј&c��p�-�%A{h���=|I����uj�:��.�T�q�f0J{ {���i�NDL��� W�yv���j�d_�E	�勧zU�d>AqbG���q@Sσ6�|�;�w��)�E�3 Uh�1Yv�̩kB��������c���ˈ�w+�<����|�C��k~�?ё�D��1[�G��vi�,!���A�A�s~E�V���`��=�}#��9�%|���gP�J���Xn��ܭ����)(sYbUWs>s��.S̾{�IS9�Uc�r0�W���Dc!E�`?Y����ʟ+���+�8��=�H\�*?�l�9ݓ�\�7')���E�ʯ̎4`�/K�XF��D'���EϠ��4 �&>�/O��!�[X�����4O	y�1�N3�yK�<�V^�qi�~^����ң�a	�ot�,�N�����s��A{�� 0Y�|�ϛĬ��XHo�18w̪������$^��XzǆD�_��t�TX���'|���B�3�~bP����EG�BA%s�x�I����#-
نEa���T�i�x����@�"�i��쳾�jD`��A����=�����KP"�gq���GD!Po_#	��)n�I��� �[V W�Q�o�Le�~�jc��� ���>���X� �9/r�ÉƢ��8�3ew���N�J��%�p{�JR ��}d�IP�n�r��+�EG�|廁Y�8�/�4EII��1`��-D��)Z5�.�(w�\�-y�-ϩoWڍ��M��وȸ��fk�xp�ǥ���Z���/g�3—�FŰ�������|H����C���Qgh�U��">N� �V��t(��vJk�N���S����V��� 9;	�dt>tm,����ӞGu�'W7:��R���5^�p���L���<�w�G�ջNj�7��r�$z�1W�+�7�^V�X�ȓh�<m�a���%��n8+BKYt��H4[�����n��	Ae �SN���.S;��/�W:�-$�lh�zGp՝D~dՀ��N ��G���0�)2<����[����a�7��s���ư��a���:u5b�p��ξ%~{�@< �Tl�(��cDJ]�X$~OŌ��)Mq����}�:����^�<�JrL��i~c�>f��b��#�@����Ѭ�>����\��s�}T�О�V�p�\�a�%x3k�S��c��w�ݜ=M����ӥ����ye6�Y���{
��Y�R��ul����8;��u2�b΄T���L��P˘%�<�D�j̈�8ޭ�1pj�ib��\��i�ի|���Rq��?~������T�3i&���gA�M�����oc�Qd�+q���ǯG�*J�#�E�{2������sWW�w�ٰ���>���=�7hc�a�Q�N��it������7�B����z86��+Ho�s
�d�}��+��]��4��J�G��J��U�P�����P�3,.E���\�*"����ד[^-���,���/�-6���T$��c��'qk���W����@j��ʍ�טwk���Q�B�?�^A��ԏԣ-��)�l}�����p�����h\\�]l|��ۇ�>����A|�_��J�^	�H)lRU��!��V݆c���4- E7����xo���+��4/k.�d�m�as?l/���p����9�e�uz3��� ��pM#U��NG��bW���my�C4_��[-^��C�����2}�ﷀ�3��^伨�n�q�U�
}jV1��,�ӴlF�g~P�J��{I��eGr�W���v�#���m>?xZ���
qV�Z*au��~��]�|D�1�6�T7ͷm�돲��  �{�P�q�D�j�!
�H.h4�WH���3'�Ss�{q����)mlS����LG��B��a�  �L~�/*�F���숄b%7���<e�\��'��e�����R�M��Y���[� ؅����jKT�Wq�H�5�o
.��$��`D]1�G ��KtP�а��z���Y�I�C�-��O����~C���1��/[�`�]1�A@��oj�����]��g�, �%M�D5�bغ�|O��g��C��7�&����h��\�#���l���V�A�"b&657��{�'W�����&U�*�OLj�-��rJ�X�Ғc<��{=p;�?�WB��u{y;��9f�ʭ�.W��Uû�O�|h?����?��H<��D�gѣ�m��dT���2����5��^α��!y�֜e��;u��@RQ�T'��ͺ'���z�<��% �Z�&Q��N_>hϧWYW���4�*>Sz��M���Y2Yſ��g:^Q�⭊�[��vٹ4[�Zl�}��2KZ�ͱ���X��w��	��}���>إlܻ�{Ua�o����&�ܓ�c`m�%��%���MZ����Z��n����Ic}�2�=<;���$K����bj%�E\_\ȧ�9���=�v
�]F�(
GI�әP���/��}�P�S�%D��u0OF%6����n؟o��=�2����Y(���)�Y��B�ts�R��#�=C�����> ��7�e��Q�q��Z�0Ě��� ����$x���� ��8�a?V�<��qo]	������؈�X��}�&�ώ~j֎;-[�)��0E� *��˪n+�S��k���ϧ(�N �7��]���lQ���+�w���j��K��&��{�|[3�y��x��?3-�s�R%���A���;��;g�Pl���}�Q`9:���i��/n6��:��	��8�K�dP&�#o�3���tR�^���ơR;rb BbY�fǎ��C=މ��j���/}�9�&���5�`�/��ϫfJ�M��R`^ ZB�u�MP��t0#xH�$�B]��	�X�'=��z�}��wU�o�V�iM_<&�^K�I: �k��r�=��u��Ȑ�_G�Y�+�]y�:]}����v�u6v(�$o�aݵ�a�m�������o��o�*c��0��Vj�4�hOQOY�ؔx�4P��:����ǩ
*�uz�j�{Ju� !�Y�H�"ny "��RQ��U9Uc����G��v0o��q�-}?Т�`\�Z�^��U��ӷ�8���h�����.�$Z��g�=���^�&�Y��Lt?�g)S�̰���@y8	>�~��"p�7�[�ح�i��xX��U�Y\� i��
�>K��
��J�����髜���PN����FN��-dFIGHRDe�5�^#��ND 	����3�܏QK.)���I1�����IQ�V��6�d:����1,��/�G�M��g`�ḉ��f���D�Hw�_|�l����z����D����U�E#��b�:�%���b�����,S;jk�5ʹϼ-]Ґ�H/�v��ۻ����S�`�߹T}�_���F����_f��L|��a�^��l�\v�W�%~����-k���SL\��+�g�'W��d�|�d~��1ɮ�Y��S[^���,�7@ ��]a��o����;0�D�<9�z�8�Bg<�fy�`R����b~SK��Jg�>�<HG�*��Z�Ȑp8{����;>��ye۲Cux++{J��!�$tM�2���ܿa��m?A��!=���������pR�4��Fh=Q�?b��#�A�ɜ��UvӶ�H.���u/�P�1ƕ���@�ջN�B��/�{u�����T(þ�%��a�r�p���G�pa�4�<�q���͋<̨,����� ��WX�M&?��2r���C���}�~7�FI�z� ����#%j5)Z��� i��"�T8م��Wc�����QN�"�,��ԉ
��Vk�V,4=0S�ڏ�LoԘ�N��=�n��.?sj���UL��E�Ŋ���d��s&���qÏؐw}|ЩV�iޠ-9�E$�\F��g%��WF^��TE�'��>ϙ�x��Zc��F��WIOH�m)�O��mGl8��]M�nܯ{c�fv�_������Z9�LPJ()�j�'��n���ڪ�-�aܠv	�u�i �V���X:��oں��"����P�ת�>�X�zn�Q��R��-wo����B�_�=��eH/!�5��s5v-@��=-�8?2�����'D�(�؜�D��[~�F�FT\z�0�L�0��t��R᜻5���c���/,	 ̞��Z���}6Gf 
|���,�\�w�bX�4L@qfd�m(��w��A=T�����x�4�y���ݗ���Y��ch=�]zIQV bI���^�]�m�b��B�"!V��#���E�4xzc�n	��l���Sy|�i��sS����h�d�%`�OZX�q+�K��c����r��%����i���6baj�0��b�×�Xƅ
'(+�=�YQl�%�[<�q`Y1�?�b�b���4��
=���e��Mh��@��$�����-%Z�!��UJ��t��P�K�.r�hD&Rx�9<A4�}lo;����7U�S��X�.-�i���E�A@�;����y��|$�	|WT�RT�oIo�pܰ�)@(/�;��Wb���rK���h�EIO��|�����&��ȭDͬ`,*��ۦ��~v��[6���C��\�W�m�i.����KTR9P2��:�b�ڑ�JR�#���������@a�`����\;�_�h�*�w#=�2�Z7o�ώ�H��G��f�z�8��Tܖ!�P�zxMŮ�o
Tk�e&��%.���b����l����9�m�zIʹ��쌞Z����<~��S
;��(�@�!J�}eUS�ۖ��,2d/o�߈�[9ؾMz�L�eh&6���2Tj�{�U���V�&c�[:��c�Nۀ��Y�dyE>����������A�ϳ"�M�2}v��vP�0N�������zyUs��YS�F���-����������v�4���܏����W�Q��7���޻Ĺ*�8\?ȏf���֒�.��-v�H��ג��/ߺ�I �⳰�����
>�`�
��3�U*�B v�Y�0Y5�^dy��� ;�3�GWǁ��_��e3J�H���������O/)mSQ�W�c�f}&�&�I1���+9��ɴ�BQh�Zy��50�P�8N��ㅪ\@K�����6��ϩOlt�mӳ��]*�,�W<�ۃE�_ކH=��I���H����pK�[�I�1�*�n �Ϧ��vq�j������[�ݚ�tn�i�<g��)i�p7�;?@o&`P������*n\eޚ6IZ,��o�o�>�cp�����@�d�@�� ���hT�қ�Z����\?UA�7y[uN���JX\=������A7��	M�u'���+�"�)���]����
mڹ��̱:�e����j���u�߻Z�('*�<������3rn�����j��0F6n�Y�h���S�|'���gc���~���yS2��]VH��O�u�j>3b(ȥf�jr.�|T3�?�g�-��5�"��S�-�5�ِ�[uۨh�(ʋ�*twux�.�Ē'Di�����l��t��5���(�ZE��S�5�uw+|�L��jT=&�N�%J9�Ic�$���/�uL/�����jl��n�e�0XƎ�ݡ�'p<F��.��;��';}YGzR�/l&B�(AĨ�� S���[g=� 4#� ,�OH)����o�	�+.��^�YX�<�I�{u���=��%���[q(��T� 3l
��V�OX�h�H9��7F��A	��yL�H��_F��Y��hZ������③¿��xf!U�����p������}��I�窽3�iv	$%@�d+g��x5ϷRK��<lQ�`�a����i�l�����Q��5�
O��{��O�yS�8�-���vq$��*�]���<
������7�C��umc��a�g�q��K���0��@�a&d)氹���1ISNE��o�*�`�г/�u�I��(�����s����n1E��z_]�W(7V��n�tLW[�ce�Џ�[�۬vUb�v��f�Ո�e���n[��;���pN׽B,��	7��P�a6���#i�tz��C��{�tި�R=/�kM�R�qG�XoEyߓA��q2\��Eq���ѵB�J���WQ}��Lh`����h3����[�l�ΰY.��I�y�"��D�ќm���i��47T@�M"}���`@���(p����m�˪��M��6%s��+S.)�F���1ai�N�����1�k��0B���H���ir*��]��U�E@�H]���%S�t4�.�l �(�~���qt8n�q�{cC�s���g���	��Ȅ����Q 
��ι*�ɰ�;��5�&o��O�q��/]�	��R���mlͩt�`����io����;��i�Ш�y��^}E���� $�ڑ���k��1E�کE_�9K��Gs�����c�@ה�o��ά![_���+6͵= N�T	v�r�;�	�R��)e�vsR�H��[��x�d{�h�h�����[6ɤ�O�2�B�~V=F�����^0J���_�F����z������B�Ԯ=�-�B��=����U5a�a�O3�G}pp
`�ղOv*9jM�O�%���r�j���io��v2�C�Ի�}e��e7{��@�F��VGԩ��
����볻����8'�6��ZC�l]ۋ�~h�%=��!R��{��k�s{���X9қ�EE�D�����0���C�q��Io�x�jnYH���>�3�*�XX��%ǈ�G �X������_��X��m��b���=י�W=��������oe:��#R�Nr��~b��{Jv�/^N�ن౔�I������KX�����e�,O(T��P���4�i��oPRQ~����7�Y�]K%?f��ӸDv!��{x����XD�uF�{�[��,�OK��%Ē�ו#(�xH/���s�\����ӭ�bB!�0�Pay姝i���t��z�L���_��yp(�a��*��h�3��t��m{Z�?�3p�貾�66�`xK�-)4M�.i�9u�[2��hZ���k�=���ۻ�b��&�wf�[���2��IX>��h�2���=��M�xGJyt����RI"\��3L���\� �m����X�[Vp��4�FS���dXt>��f>�}>G�c�$d�䉦�I��וi\�.���;z��/��rųEK�:j�ٟfh����qz��9��z��B�&��5.�l��pao�lY�J�F�1f�8<m M�l@F�k�$�c�zP�`��X�so��FD������3�g�~@"�l:E����O�rw�=��9Ȱi�LTǒ�l�����O�v�0TH��>��V�vS�z�+5N���*e�	������0�tM�_�1 ���cC' x6:&|Q��g�h��| ��6��A�'�9�Ǯ��vy���yBO]M l��.�^�S�����_|�ps+j�G���g�����%S��Z�e-Bo�1g�w��!��q=�`g(���U��#�"�bV��6�	�� �v����e�'m�=����D�GEy�	�I�3��q���Τ�x�>��[KX�!�`)$������-y[S�'��l�y;M{�pS��u}�ɷu.EVe�'���^�7
R>�
�Ŧ�/�����S�ߥ>$���`kL����b���t��M����
�U�J�jitD/#��j鏢P�����d��:���\��4�nx�h�c'�i�q`7~Q(ˤ���}��h������@?	ɿ=�םۣ?����X#zx�x��Jͷ�>t�<�O�S��Ugf[���ȇS��l��P���;�'��[�`��F�c$X׍�O��:ГGX�=���v@>�i��$�1'��p��f���8-����`i<��q�0m�J�^M���r&��s���N`��WU�z��t�� 0*��4�`k~B�{
cl�2೰���߿}�Q�@4y�AF�����_&��@�	ݡ7�j7�uc��қG�I�!���B�T�Y��F{�QF/����S�� R���۪����T��:C.68��V���nV��)1'��Oh��slf6�3�j��{��t�*���Z
�a�	��&��<T�ݢ��:L��cIC�ߧ�ԟ�肐�Pt�f���X�׮�,��O��Ե���i��>�r�4�� ��l^>�;�*}�\E��z�u��u���K~#���*$�ֻͽ{���ر�ϔFiM���S�����#Z�CƂ��ﯗ����0F���lB1�ƴV�����
�p02Y�Rq��n���KeQ��EJF����w����]��]HG�ejq���ر���0%���VK1r�$�Ⰲt�6����M�����h�ͣ$� ��M}�έy��;����I~�Cڡ�U�i����R`����|ytӗ��E}D�H��[�b����b�Dn��e&[���Vzǎ�ҋ�D��|L��X�Z�.e�[��!U��%_L?]�'ig��D���uVk�sc �JՐ�9���:�^X�zҳ8�-�%�yF���i�����?|�.��-�N���$�x��:�I�z�ќr�|�x:w���v��\�'"���m�A��&��>�_�^�M��=4r� ����9B�L^��~/���|����;U�O����8d��}�@w�J��!�_kuu7��D����!WAϰ���#~�dy�3���~�8�FBgb�E]��2�*��d�6��y��!@�h{��E�vK��&�<:Ն@ѵ���)������2��'^�8h9�(w�D��U��,sh
��.��8��C��D{roz��A�����A�U�_�w1��i�����}�Fw}�/d�e�P�R%�%�ҭX���`�wg������ݚ�K%(גk+�XO��]�\�̰���;G������
=o( =ln3�ng9Zo@D	[5�Z����q#�:�npߛ�����Ɔ6�s����G���m���)J�h��GE
$}�(W�Ce��j�h�ϫ�I�0��#��4[]�g�a�~�=_����$�U��6ŋ�%'W��X�p����_���^��|�t؊̞ˡ|�h�Fr�/L�؊��B�W�k�&�S*��֖ՊZ��Z�py�C�uH��8���pQ��F�qy�	��	ut��<��<V	k ��E�p0f�G����+��vU�l��gkzll���,[b�BV��^�{;�����'`��=�N	�aV����@�7���|�b�"���?|��X�v�M� ��+o1��������D�?�Rܿ�!먔F.���97%�R�@��'5%�і�t���? ��'!H�`*�++,k��������E�Ұ}l�����?��m���q@���vt���ڴ�lf!c��ߵ$AC'�dI�SqA�	5��[�#/�������x��<8�7N1�T�|����YX4bϼ��5|׶�����xx��>�U���p�(��Tϝ�!XV ��b\b8�Q����x�w3�`�D�)
�©թ��)5��1�<�	�-R|̸��w��&4��j���~����<D���Wڊڰz� 6���J��3�s�@;~I2�Wp���������8봵E^\9J�v�Q�kʢ�S0m�`}�������hD
9H���v�2�2�ж`"z'C���L��CD݅��I^�� [�?�%5�'��؛��
R�3O��,����h
_v��1�Ss�T_l�����TfJl+J��0e���X�~�5O�9c��ւ���1�=w�!L��7���󖯾���^C���g�Pl�}�?Pxd�(�̽��F����������q�1�f����)
��c�
i^Bd��Y�g�?L������x,D�3p�.ܳ�k����$�Ʊ۞��4泑5�	�D�� �_^�ɤ	�
�#$\xH������I��7��8�解�/80=OR���{��	��l���>���������u�8� ��v�aU:��⟓G�1�zx�>.������D���&ē�qц?��okF��b���J����P�����N�%h����[5�׳�\=غ�S
�3�=$�S��q�*�_����5m�`��FO�N"���ڴ�F]s,'�����qA�w���0;�|���HR��Ў�O��?C���z��äר%�'�1*��X�}�oar�Z���~�d�`���VA�!#���_������r� �X7��&$%�2c4�����p�2��
�#�L��Iw|���YP�0.�ɝa��[��ì�&�9�h ��D�1$Wc�y�� 
��eE������j1!+9p��i���W>�=5�e�z�bk�ƿ{x��v��:��>Pǹ�e��FH]�I��H3�{������c/B�wm�fd�+4�Q��)	ɠ��(%�l�i5�=2�����T���M�[��4��J�|���BC����1JVǒ6�h+���Z
�@��ސ�$�vռ��& \��3r�܅�V3�֢X@�����(�d����I���/�G�ϵ��!�D���D�z�P�����:�ywK� ����Ǜ���-��A�E����N�A��73�Ƚ�����������|�C��`2;<�~L²��K�qMt�����-�+,��"���k���'��(���~��]<�!@�`��p���(G_43!��m-g�UJ��<=1�0A�͞c��]�z���
h�&ݳ:�|j�'y"��]UYp�bZ� ��(2 7��5P0EwX3{��*��^�X<-ԑ�F�j�+"���jx�WBj_�t����+VIwGqѮm�'�:c�\�YiI��h��8j7�}��	r�,odyC]3�����!.�U����֔  �Q�sZR�J���_�Tπݷ��e)TYE%�� mo ��l̖�m#E����~�f�c�A�Cx�3��e��>^�iP�=#�K1I_��4�z��+���Z��F�F]�U���@)���f�z�Ȩ��$���
�@���P*�T�Du��|�q����=k���O�K]"@Ee3r\;�]����o��Db"����C��a���̓��VW��R]�zƇ�r�-�Ia�6�Y0vR�bq�}�PǬ��� �"�]�߰�7擷8��4%��a�.M�!⠑�ǣ��b��P���+Es�駃:�0�cF�h��k/k�Tg�vӆ�y�����#�GoE6ע�DƟ�Ym�U+n,�4T~����	@9=��dz�t��ҭ�?9� ������̶��$�b�∎�9q`�%�������+��������QT���=_o���5ȠZ���~�n�Q9��H������r�.O)Vǒ<E�l��&���s"��V[,��L��;�^�VR�$I�]����4/5T*S�dU%�] �J��|���z��&;�6~m4�������fG!8	���X���zf��$G�I��_Z��lʒs�G�/������7ӂ���@/k
�}��X���BX�d��DX)���.��˜ϋ-��h�g���B��5g�������Ǧ-�E�uO����lݚ��O}9�ؼ~R�ޥ��n`:�t;l6csA`tr"˙�����.{ms�*(��'�4O�|�oڗ6坳�Z� >��5�6v��Z�I���F66୴��̻P2�n߰T�{7�p�
G�	��{��L(�10�@����NÖ�B�:+E�U�\M������m����R)�!ͼ� �w/Rqb ]Qn� �ʍ<��LN!��N�2����2`�
o���f-(,
�|
�QӣV�*�_SE�G
�ddk���5����"�]QM�g��h�	��s����='�%]2ʗ0��AXp��/F+&����S�_!�Y�*+nk�۴X�5Ћ =����3ȷ^nR�_J�m�0�J��T�� d#� ;����b�E�z�0k�J��#�!��3���s��P8�N2�}1kф�3�H��/��2Hz�<�QX_���ĄJd��#,yt/�a#؇YS���Np�@�"������wb��œ���-ǳl�ݔԱ�]���Sy�J�j푳�1\Bx�>X� r�~#����Eڞ��6�ҍn���&������a+��v�5L�7��B�y3{�����/�/f�P�x��B���c�:���ۉ��Ǟ��ץ��X>���W2H1S�t���s��Q�wP
<5X��,y�c}]�����@2T��?5"��벐���G�?-W�%L�ZST��/1����k�J��9�dQ���K�߶Ny��5��BǕA��w��h�ۄ�iʂ4�Mh��e(/�b��c��m��R�����5���%Q+k�i��G�!�ͷ�_�)��8|+��V�B���O�h�c^5���"1�|��z�b|���6t?��,���R�=% �.���qb�ӻ�Ǟ[�b)Y��htO_�&����)C�&�X`k��Z��%'��~�vyl��$��vA׻To5%��*���Ch�J��� |�6Vr!N���#�v��9~b�:fqW�k�J+1a��}�zMVy)M&]��L?�iT0��rR`)��䩭QY{���㞊��b�*`^��c^Wi ����fe�Uj� �͌>p��a⸛�t3�����޷la��ݚfo�W9棐w� % TZ߽��G�Iɲ�x����=��V���{��8N���?<�R={��>��޽��v:������q7�q��?U��$�����Z��_ە����y��uUc��5q�p�S���TCA���\7O]���k���)�����\�tŇr�(�Z�(]��Iʺ}蠊C?���:RD�1��$}������-������T�@1��A����+K.��w.�7l<4:�8��U�&�e7�(S�xU��b����N׽d��n.��*G՜���Č�܎j	��3V�5v�COIu�L���|�M��i�0��� P��h��$$
A2~�����"V�2�b"bR��`W����������p�^VRå��;$_MR�v�-�Z�P�F�&�C�}c��7���^ӫ;8)�[y���w����@�#�j>��}��������eJ?�r��n��[&{u5��G[�DC�l2Y$.Oq�!�����&�c:lW6��7�4�S`��|�	O����nm/��a@|������0�/�8uLG�>򥯑��<6bDweO�f0�)=	��P+?7�W)��; �/�
�(M�3�B����ئ���0��?<4/P)�����O���	���ag�)6���	�Gp�z��#����o��f�:l=f����`O�(/8���9N��i'1!��z�c\\�+j�ȣߧ7gF��%�/�gĉ����W��p�ܭ���9���a���m}桉� "��K�ǘ�I�S�R	N�8#�S�}O�By����a�@xړb�8�`K�}I�����cz,���o_֞��B�g5�Sd��~�c�<��3�7�(J?��_:�h�ʱ���`�����*�T�I�hڥ�A4���[D�C�(�|�:�}i#5���=���0G���`�ħ��?�Kړsi ���Ov�p�>��㣖V���� c[���b6#�� �=��EhR���wgM��y��p��%��B��ǦC���7��푾�9@F�u�VC\8gO��ر��.#���	�P���� ����1p]Э�Qw��tʎkQG�}�1�,l��Y��ͼ�0��dNEL�Ogj��B;���͹=�#g���૾�G����N�Ҕ}숥" ԘK{�PH�M�u[�o�Yݣs�G�����R�R%��U@��5��H�R�{�(�6%|V)v���'q�o�H;C�U�-X�|��&Ub���8���4�bQ��e"�ؿĺC(R�"�x�W���+)�Ey���)����ؔ��X7�5��;PG{[8(�N.
��V�w���*�׻�f�
�a�9^�@�"��rz@��rK��R��r��o�P�xW�=>WF��d����cCJS�Z���$�u{���f�-L4K=����Ӆ�z��tn�<T�"9l/݆_.2����.���@�"x��2=�����n\���Q��h� ,;1��l��2��x�@�0O'aGG���|�t���SD?�`�$.s�3=aZf׸Nz��<���5kNj}��ҹ��2�,YD#�i�MBF����?4�1hN�4F)!�y�}n��Ȑx~&�
֤MB1*(���25Y��m���Ԏ��@�Xϰ(E=\q���{Vj=K�uZ��g2����Rv?�s�U:$U��<�zN�@�\	�t�������j���"�D�{���;f��L	TF�*��(c���*^ޞ����V@�6ǡ�N��%�Y#�@�¦;�s�9�/�[Iv��3�3s@��+�X6s���g����T<y�&��e��B?�e���Y&#�mf���s�U���>g�	�ڃ=C�=&�aYK��А�Zx���&�T
`�c8���uv$��?��,X'�"���ـ�>؆�ӟo��ʶIR`���%2�Ŋ�{zM�(7�2A��rM����A�r����������ʹ��~�5ф}w�2;ݮTNV_;���5#�Z�'s�2L���E�GV�Y�,c9Z�)}S�xR�2&YlO����_��e)єvh�dˏv,�cH�e�Ad+w�M3�uN�!#S�Y5��/QZq}ֳ&�=-��g�J�X�\���{>�X�#j!��
�E[�,��AYb�%:Q�V�;1~aqL��ڛ0��6��wHnPє)�գ�� �6^���$v\��_��u [^ʅM���h��zEI&�#zWB	��}���)��x�z�\��?ƚ\4-�B�p�j�5�M�GZFC
�|���}�=P˔A�n���r�SP���4 q�n�F���	��Eh�6eIOf�q��d?�9���������<�q3�cԏ4�Jn4�]���H��f��m�i؎���h�����F�y�_jgŘ��sS6�N7��XD,Q��3�.�|,�KݗL��^�f
��hPz�p�Y��ud��,�x�[c6}����kTJVդo i�:�j�<�F���IQ�F�l��I��?�G0��}��&�Wj����
�p��'�t ��	j�e�1��n���n!�����g��'K�8�2����~��y��%���/ �)ʄ�}��-o���� ����_�	�֤�h�WPb(�ᙧ�v,�YcK�S	�e����!P-E;F�J�=�us�o��2K��q����3�s,��gt�����j)���L�DFK��i�+����8�T&#�d[E�fVj�]L�&�V@���;��L����[*�#�m��t��akw6���s�2b����&��a��)�H�x5 �0F�~8z�z]��tW��7;\0e2��x0�_Ғ�� �5�����ζ#_��~��8�>ko�/����/(�cfȰ�4�*r���O|��*���p��=�v���O���l�h
�8�u'�\�<Gs�����]��N�@��M��AB�5�3NM�ՎJ�YDa����R5�7,����Ղ=Y���� u�RPz�����Ue?����aK�����l� {"�&�e�T���wF��\�7���kR����A��;�D7˶��&��/a&Ÿ���fH�p��k����A�Q�ސ./K�8ƥ�}�S�� >�vR���b"u�2��*UYQC�裪�߰�x9V��W,�P��6tIwv���ђ��B�D#ϛ��a_w	7�G'���ă �ɔJ�{���g�/�#pZUb���m?����"�{���m�/�h"^�0CI�T$ɅЎ{�rʔ0�/��+Oz�0������zS�.�a��zH�+��\�c5�ra���+ ����R�-�p���"&���$a"nA?��l��`�i�>^�{�z7���Zb/��p�OC�����I��v��ΥwZO8�\�%#�I���I��<�χc��w(��i( ,�X/5!�'��*Ɵ�L|]�|���;��ۧ6"q52�CB�~��\�3���B �?�:]e��N��_�	^�*.�ۇ"5����B^(
����n����T=q��b��`���)�@��7��8�SF[�W����3����,ā�cޖ�vP}����/�]nb�H�svo�v�z�L�$��\�cc�1��*�z��n0���Y�TB=���j�ÀY!\Ť��w���{Q^��ts��x�(ܺ;/��e�M핽=�09�"�T;9�ԇz�,�8���t7�M�ŕv�� (�Qr�M���r5�j?DH���}���p�:p{��#:�_.c��A�s��G\��Fd}l�en3�?��f�\�S�Ro�G&�sfW��a>}�T���\�<W85�.Ҹ�(�  �+Ϳ�����t��4SG�ƞ�S�-aK�Ȳ@�%�|#�~ ����'	�͞����m#ޠF�$�1�)"�
��M8�x�C�����,ͪ�z�8re�
�1j�$ы�Xsk� �3)��B��~��֚t�Y�(�U��Lݶ�c�
� ��7��{� u�[w�Mr��an̛'$y@Ih+㏫ԙ�OOלV���:��m�������<�%��Q3���#�Al����Z��B�0��"��t���m�"�~�i�G{��2��)�ݗ�[�uCV�w(�x>�[��ȃ��̑���Y9���yx,R��uP�$�G�6��u�5�H�:�Y\������כ��"� Xpp%"�~n9�@�"���q[���q;ߔ�D���g�i��r���V�%����a��d]o�����Y��V-�=v�����O����	�"�/�$�R��߻�xH9�]�q+���f�����Ք�����6��TpdA8���TG���|��%� QmWA�J�ϱʨv��^;ܭ��G	�Ƹ�:�.���S]�o1����䄕r�m'�4��:*k��-� OÄX��L�B�Ԕf��Vƥ�4�������5j>�P���ߊ���iJ>�uw2�~>e�� 2���ENd.+b��J�S�B�"Ϗʄ� B�ay ��Q�A*!iIؒXv0;�R�~�](��;���#PG�\
�\pH5��t��!R�^ּ�E��H�����ǀ������Sc -~�h�Z�8��f�K�k�!�\��ۛ�	��.l}��*�P7���U�0Al�s�e�bdlo�Y�Ȯ�R�#�-!�U�9/x��ġ�;���ڣ�B���� !��%�Jh�PF��y�2�*����0TC1��F��_��y���lг ��֖��S��T�B�����xh��an]��A�w"�4R��7x��l/}��G�!Dۑ~��Q\qF��������cb�H5�}8C��s	U�P|'**�?�9zYfBr����i��V �If_ �L���sڶ�YǦ�-L��K��q�6�^k�#
�Όe+΄����Ѯ7 �B'�a����B
a���l�B��ckC���U�X�K��;$��4�AU�\��b��jY��Ĝ:�6�A x�d%�q���|���|�K���,�W�A^k��;��r���Bڧ?��%Ce_�<�|ъ������:��*L{�$�c�.u5��!�Y�&��}BYv��|���%b�l�}MYC�teiL5�s�R++-�j�Zk䅔�4��׼�s��V�*��=_[w^.STV�.���"x�f?)�?�C��(t@Pzw�7�o"5:e�F��i�oSZUF9]ċ����)kfǅ9���D�b<SAŨ�����a+��,~LG�pO�QXȭ��Mۚ=|��1�����O�,6�f	hZ#�?�������_;����]π�Ƌ*S o�#�!��JC5�^�awf4~��n6�-f�k9j�c�7��UE`r"��I|@�C4l�'X��	}�Pl���᭲�{�0�U����fS��$ ߅E] @Ѯ��&�1�~�C�^�V�I/�%���U~��ǎ��]b�m:=�{Ǒ����qi�76�����_�S�.�M�{J��WM��8��e�١���6��:���p��6�5��S�_�ֶ��6B:Ж������J}'ix�02���ڜgIq@�����*|b?��yE|���Z%���Gc���.�S�
���e���
%��B����:3���X`O�[��\�<z���G�)�q�cC`CG0��Ǉp�AY=�):$ [:<��}z�o[��q_|4HuԜ�@��W��'�5���؟ETHR��Q�������-e�v>���Ϲ��by�C����� +Pi���D�q����b�u�$�U�9q5Z�g�ʐ[��`��t��#��Le�������G��IRS���K�Z��?�
��QCv�!��?i���ǻST�hcOR���Z`�)�u�`���rU������d����B"�M�Y$mX;�%�)u"�8U�}�D�OGZ��D����fk������i�{�@B;��e�H���9?;��s��Q�5���A����C��f�i5x�'�ܢ��S�FxZ<�R�����v��\��a����I���3�p���҂��Ո��uMC|������RFi�\/�?�B�0'cX�٦����I�lol�e��п/�2�6Fí��FB�+P���.	�?$6��Po������	��r�;��+$䥽u<�J��.;��G��Ӄ �\7���P�sګ�~Y�c��@2��'wwu�����=L`q�R�͝q����$��߽�����^���I�u� 7\%f�p�����o&$�Wi�e��B.�t�ܺC�?�uUg����#C�K%yyU(��E�R@�<�-v#������8e~��Z�����qİ�� 
�nG�R�m}zU�`�j��I���V*�#���ϰ��"<S��E�%�D ?���}���6���3	[����T�|��a�/�
���G�&ILd�(�i�XOectj���X��daد��u)nZ������1c��ZFn�#��(o��l���e�N!A�}.�L�`��n%f\����������yE,�rH�H� ���e�&4C�1jU5�5r���	p���[9�m���#�"/OY`����2V�ӄ��d�T��x1&�����7}1-�.tE��Q��ӿY)�1��J�^d�C��Ҥkà�#�q��,23(1.H0�͉���l_{-IO{��8�̓a���Ҍ�rf�#�Q������[Yv4���,�.�����RL�v�"������b=�M�x���[�I��Y,���D	����!�E��C8$ǆݔ��۹�Ȁ��x῭c0��|�5)�(�~b��44��*��l�x��u��0Յ�"�����ڔE�(:z�!���k)�����?h�R6
���_2��gS�&&/7�w�Z�3�X��0sv*<R�.�E����M\��v�� Cf<�&�h��a��sG\t0z5�&��7�ņ#]�_�r	�;T�[d2R۝-N��P델�?A��Y�!K�\.ud�Pk�B���ֈ�7/6���f�2���p�^�N�VP��y��|�N]�J04Eؿ�mͱ/������CɴO�g������'��ⷞ}@�4��3��ig1������l����`'P��~@�c�IZ��P���8֎`;nRY�p�C�AnC$����e����$y2��
�H>]W�ٹ%y�����``�A/F��#���o�t�*��5�Y�>u���Ժ=֓A�}'p�L�V��H�¡�R�K��@l��5��}M�rӣE�S�~#!��A�		QM�SC��МMB?U�in-W�Ck�@��B+�W��k�m /aY�����3�@����p����J���c����ö�����#��"p����G�G܈�	K���� ��oaN7�j8���F��JA���j�Ӗ�춲[���/B�io4{�^�M��^@N�o��'�y��g~�Y��Í��O���.�@�݇�*����q
#�4b��J$�D F��J�?V
��(������+����̓4��>��������E��X�0�N�J�dU>�@�l�G�,�N	�{�/㢞ˀ�=bNK9Kxw%�l*hƪ�o����`	�u�;�&�MF�W���x-,s��1�4��P�)1H�▷�V�V�A0��� b��ۚ�q��'���|�81�.��G�&RF��q(1�Q4U����a���2�k���RnN��[��a(���}f���� g��Z�t@G��:Lߥ�Z ��F��rg>����X�2DCu�-3� �(p�����}���$G��G�Y�"'������;�CI`��ď��D0T���j�_�����2n##<$���PR+�����PO0�WO��H�ɴrm:�2_�qUC��=~Q�K�e�|��F���ґ�ꝁ�|sOV�8���Ds�o��ڡUdt�M�j�S�f�4�
��h3f�~N=�$���%�K;}h'�����W�5u.Ƥ��V.���u���M�)#��F��O���dߐ�a����6��~j9�;K,���s 3k�#���B�Լv��&�*/�8�Tl���c��	6��wsXm�CV3�w��P�p���{�E�#J�콛]��1IS�T�� ����o�OO��$��_W�o��z�+�.�s�N����F��,��>%B���=������AlZG�*�B�~'�(:P��A2����JY���Ȑ}�f���:��7�Psl�tSo��&fJ[����c�T���-�����'�2(Qh�fO~�R\{.w���>
pp��LN��Eӏ�vw�׊�tm�����6CLŷ'=Q����B/�T����>������wL}Hʮi�y��?9��x��U�ª|���eǞ�~0�b5g��7ϹGu�U����KD|����{q������zl{��_���'2���ԈA�$͍��8�T�'����AF�ֽ�7���.��@1;W]��(�"2��V;,���p��uH>־q����5凞�*�X�J	v���c��\y�E[�Xw��#a�~d���_�}��o �'�xh�[&}S홽�&:/�#6h>c7w_Ւ��+*� �����;:�5���A�Z��V���@:�/��S\�>T�㛼�!fw]�w��NL���&v���B�7�R&U�xIB�<�A�涌6�����~�僀���m��?�
�>�{�FQ��J�?	gx��>秥-^Z%�M+Х+9�)uo��X���ո�:Oy�[�|]���n<��IVh��AY��5]����X�ˆQ��)c���d.*d�=ׂ=�߅L[/D���:`�kTYbBX��H�S�1�O�/������ⅳG_NUo� �U5�*�u'�0����Ap�����4�!��.Av�0�R@MJ�64:!�ѡ�ֈlp�cœ�D��46��CD�Hq�b=eƺ���̪l�J�V~jЇ��}~k��P��p���� H<k�]hM�P ��?}`���
�.k�N?��7��QS9G]]�؁d��(=�E��?&M4<c�D����>��.�w�͛F�Kc�����iU�X�2
��T�h>��^�8&k��kn%���p���$%2�Uw(�&�T��l:A��2�x
���3�"' {�Í��c�MXl}@ī�͉qy�g^O��Ӷ���q.6s��XeY�X����A���*�V�ֱB�M$����!�Y�I�?�l����i@�g���c��烁�J�F�=��
>���<���bU6�0���>6ݜ�'m'5��_sBgu��l�a�H�djѪ# ���|;��vA�ό�/�Nf;�p�M}$�\=��Q�*��c�����~̲py���ґ��Qx�j�e˽Q�Є�"3;~>3�=!@A�#3Ё%��-�_𒄟	���-�2v��
���'�O16^���˚p�����jW�����NZ)��/�������p���m#u�ve���9��CN*d�Y
ƯS+t$3��aG����]�O�g��`0�*|�D�nʎ�>E���z7�i�A!U����*Vt�ҵ������ב�/]$1��8/u��4Iº����NR�m�_��O��"���H���)p���z=A�]��i�i,�<�yX�NSh|ku�d���DU���B ����t�--T�4�Ù0HEB��V��)fD�����uI����k��Λb9b+e�DnI�gk�O�IC����h}�=Ä��ܽ��y�?3�ut7(F����c���!��xaZ�~͜����Ԇ��%Frk"���=_�:?2�b�wU+"Ы��`A���1�ym}�bfk_�_)dp�~zw���w��]U�Q��$%� �B&?�q��>�y�|iW_�4ZH��F�֟��f���S�1�!�)a/`�n��9��j�Ou����6༰�;���/��^.���Y�&RT�o��E�@��OKc�}�<�oA�E���,�H���A�p��~��)�����9o��x[W�ێn��9�͢\ڃW����zd�Lv�����r�����>Eg;���rk_�m��C�?��9k��Zp=�U��1!�h�h�G� �2�I�r���U�:l���3���n|�ad@�g�t9G�9T�j.�q�G_���}ĺcr6)�rY�� 9�nM� �!D]fcC�H�Ȝw�<2�@��KΡ�>�|#db�(�䮖+ْ5r�.׼�A?	\2�A�ԡ�Jbj'����w|���G��?!�ip
�A?ǖT����E~j�k��L[��b>�؃�������+_�e�W2զ����]�X0a�����q5p
�r2DD��^�d"�*3�]D��rZ賤t	W�mM@Q��&�:�N�����Q\`��5p�#r�N�����ū�Ñ3zѩ!Q��pol#�Ϭ/xT|^D��7,h$�b��sZ��^Z��gJ�~Jb�硗woti��YJ�h��t�n)���udB~ҁ
'��:>"EKlD��j*R��TA"Jh�eY5�r+nXy��X�3�u�a�q������Fq鉜4�;mf���zm�}�0�k^rSY��Yp����p��N}d(�LP
<r$�v�q\&�	�8���zJ�/������:!���2{V߃�������_&x��ɕ�x`58솺JN���J��H"��Vv��'����!���R�2�`�, U �����ܼ���
|u��T��p�rM��uZa�5!X�A�����h��7J�RE��R������k"E�)k��O�ݹ*����G'�V��z8���b��Y�����x~D���k�u�吞�?�Fu��8�� �rNJ����]`�g�y��s��d��=wmg���3�hY[��,�f��y=֕�dxݪ#�[�J�o7P���r#s����m}ƭ�u��	�Z�j�-F'����M}�֌�1�&r�LA����d�R�,!ؘu�:�mk�>��p�!��]��^�W�{e�OK4H�4-�eV�=�g/O���/ζ%��Ԁ��ظ�qO�Ǖ��W]�����Tgw۸��m�{��ç�u�Jv��F��.��d-�<�o��q����K��ό��)ȍ��Y��z�f��t�c��S�'����B_��e#;0,���A(���Q�������� �W��*�/}hY��p�Za��q4��Y�J3��3�$����⛺(I�6�]�A]���7����蓺�@dAlYt�+�n���;)�y��jO�����Ԑ��'̅ouˣ�+y�W�C�Z��(v���Z���V�=��N%�e%��!n��H���^(�_�w#���Eg>��:^|YJB��q<1i��Q��Iݎ8OC����S�x.���[���P���L�D�f4P6�%{���gp�ʻy��?t�)*�UDQZ{�i��|
�·#	~?;�J,Ehޅ�K�����r���y�{L���Z�@��+�?�����������<�f�OC"�9�S��K���B��#������V�nF �Yz��%�eZ�L�B�r_ץ1tR�z]@~g�W<EL�G�^��or�*��gN�ύ�q<n}f�2���r�58��Eg�a�ߡ��ސx�h�-42;�!4z�%��z�A-�d�M����+؎G�Ǵm�ۈ_k+���&U+ey�+:��x��w؋�u � HC�=j>�xL|=����B#e�o�����rB�ƾ��,x"�4#�bΡ�	����,����z�ќH���WP>�/!7��`��Lm�����.�������iZV��/ҟ�4j��V*`H� p!~� i��R�S�����)�2i@�����}�g��I`�F+F�:�A�;�D���Gr�����m�"�[@�U<n{���ɏ�)}��-l�rn�^�\�A|�Irf�vn���N�S��j)=��?|�����`�XC��mg4e����g�A�<H9{�;���tώ֊���VL�X������\~�0Sr��D�w`��3�gO~�H�9E��:ǈ��;���E���~���&��+���s������NO_b\[���9+_4��*I@���2T"��9�#�Mt��� y�DO��y�ġ�N��:�X��ų�g]��-l�D�^	e�A�+�l��y���Z�p��v�q�cPv�����[���c�)lq�v�j����4�QU۠$��^�w#{Ҿl[��K15X�m�eo�Dޛ��s�����oŝ]Jԡw�J�P���]��[���kM�����$���N��Ý��R0��5كm�lS�w��a�2��R� ����Y�|�&����;<N�����-�&���4^�>��La��i����imԲ��fS4�Ɂ�f��>mҹ������T\~,�j�s�w��n��Jg��C`*(�B���z;�$���c�x�e<^^I}���x�c|m��%'S0�iw��[xPB�������`d���T�7�L�c�έ5��oa�i�[5�*a�\��]��0�ۼ��ڣ%�/��9:������@�����Dd��䑶�n�Xk������6�Y�͊\����Òj�j�P5Q�7�O��Q6%dͫj��IhT���6�6�m,'�����X1{�mϮ�Q��'�w	kN��٨x��邇FG͆�s�{�n
,s$'��_�;A��2׭� �P���� d��*�Ƃ�KJH�A4����O����<�i&�ɊT��ؒ#���-H�l��;�A�O�|O�����8��";�����űwT�t�������<���vl]��؞�)
����*I�ͰTY�����
�b�#
��Pox۾��w���/±A���O�s:����/_��󆳒6���@:�K)&���~�[g� m@PT���� |��)O,���h/����>�ˆ))���tܐT�F��_/,oĦ��zh��Ƽ�8��zZd���n,��ӤU�5h���?���^�ʣ����M����{; ���I$<ΤH����Ȉ�qU�M�#���ѳ�����A�w������|��E����k�Q�,�H��5Z�C�%>b75����&6�%�ry�.Z��U���/ZI�lK�\t��z����Ԣ�i�U��-9��d-W��!)DJrk�!m�MZF���_|e���X�����/0LIЇ����`�:{9�N�L^[�f�]�(2I�����@�;R�Ϙ��v�QB2Д��$�e�#��;d{-�f�LԔq�)�0������t1��M���zӵ��0%P�j}
��;y�h���Ѓ��r�sXe� j�,5������S�)��yIJ-� �B3}���G0�W# ?���c�!�bl��ܣK-����r�:K�/�S�\>,��������&�ӟ�<�f��b�W�O����Z&�H������<PC�i�/�6�h��'l>S���+v��F���V�B�� MJf��[C�k6�
eo�zD�C��� �
��W�2s��|�9x��h�l��1(��ٗf+a�D��yF ���,�I���FCk	����	���%��rSJ��z�N4_�Nd1�����F0':�ql�Fs��F_b��b��\
HޅQ.��_)�O�\+��k������2k�2g�ZVp����6*{Z�n�D�Y�!NS��jT�L8Bx��ݗ���ƕpǇ)@���,�JPǢ.�Vl������f��C��H�v�Z���}3�tq����<Xղ�Gv:���I#��fy�7��d�6Vꣽm�̍�U2��$|���J�d�o�ee��z��Q7�<�ks�m�R*��su-�e~i��#}��'A��[�VB	�l]M{�g�����٠�<пk��ۈ�P􋳧�k�H>,�m�
	��d�� ��?ޗ FOZ�?�fki)���dm��~�
�ۊ��9����P��,�(�ƛ,x������
��ed#�K5���M9E۪,,�3����%��ե���J�5JqnA�b�`�_q15�m�ш�خ��o"�Fl�~�
\nཀO��@;��*ʛr�٦\���z�g�@�P����Ŗ]��D�n)U�|��gO����b�+�K��O�ڕ��W�$�Ud��*�*��Kq�6`����հG��o&�D��Ǘ�(:�H��q�,�'�R����2�Ў��mF��7��Z�MZ�ؓ�=�(��o�4n�i-[e3�7*ڿT}'�Fb�1?��t�^}�_����6�Щ����41���@�V���o�&�
/�C�y5?L#I�ⲹ�c)HZ��ni`�p���V�3�3��Πx��YX�����d���q.�5�0�~�ʹ�rb�q$�ta�^8�k ?�*����NT��/y�2���]h�؂I�`�2[�R���#$c֘)0*[���+�����0�C�V>Y�2�h�Za��8��;�����t�)��|�e�������킶;Vf7��/\�t����ja�j1�"e��_����"ﯲM���{�~H0����e)͜�
�S�F���..�<eWܣ���^�F�n�8�*ΥY Ns���OA�n����^$�^ꐃ�Ą�: �1�mi�C.5�sY ����lBQ$��X���.��y�J���^�������b(R>�Bn~׳�4�����'"�j�YnSo��Ҏ\�Q&h��ݷ �\���k>���U�2~lS"��y�q] �r�Ga�/�2K���������H5����)r�5���ۢ���[>��1^g�$�0��z�Ux�x�>�S�(�='�ح�̝0 �p\X�:�֍L`]Gሓ����R���������r� �3ŅN��7:�4�E�,̖0Oȭ�;�4;,,9} ��L��Jrg��x�+#	���mS��\x���艛3�Z����؀؜�~6>9.��X m�l�*a����%�`�DS�J����;`�
��՛�H+k���gU� ?eMRS��b�84��.�k({r ������z�ςh��I�g���%R3_p��7	J��Q�C�)���	(�����f�*�>i�����iJ�e�K
�����ZJ[�`6C5�o�b�S?����ӗ�sfl]�ʣF1�"���ہ�UP��<n
�]�L`�|*=#��z�ף�h����5r�BFʆ�~#�?����#�؃w�N*��Ɋ��U�����=ǪdӆI:h	�I:ٶ��]ȥ9]O[I���w}Nc��f]U����n���B��8�9D:В?`����5`6�"92-{�]��ߨ��*(���c:�5s��?�Fy^����nA��m���ݪ  *�wg��}p,�'�j�3C�:ltll�M`�I:7;�0��O��#�����o�!�o�[(l���N�T��!n����#e��郵"폶�jP���yg�lk���֤  X��+}��3dbc�3�Q����T�*ey���SG.�'Cӵ��9T���$#�Y�u�\��E ?��r{z�.�a�Ɗ�`���V��^��3��,����l�8�1�[���lO�*�����t�g�r�Ɨ�'� �+k;�	���ѧ�������P Z8Wi����A��ҭ�{	�]�c�
���$��7�:7�<�y��[L�� ^M�m!�iG(����؍]�{������ ���B��	�#�^�[(�·p}������WA���@�Z�?xĐcy�e/����n���G��B���5L�C�F�V_�?B0�iN��T�|psZ��Z��qK��J�@t�8�dK$��,4�6u/�������߇�Żcb��D�B����Wh�T�3��;1��] ɴFp���qD��n��S9O��/�Istz�WP��|�*>A��H[pg!uH�]Bm�MfB�#+'-!"~p�Sz�m����D.Y\�5q%�V'��։,��Ɛjm*!�Y�@����C��",�:��� �w-�M��<p��3�	�[������R�w�KE���;�]�RY�);=87��7K�~�֩�n"[Nk���&y�Ǡ�q�&��jPǩtS��a֖�/���k��qwh�h<R&�P��`�e�U0�<"q`��� �l����k\o��I����,��G�)�y\�9L���+9�@k�]i��WF	yF�a��
����K�],zr���u���2�cݠ��_j�]�ٕY��߶ƪ�~���AG?&ݹi���U'��X��n۪(ҭ�X�s��%p��xV;S��ɜ1zvq�[�%�#��Ь�5.��T���Ǟ�G�0�"���D��/]���~*Z�D?���U��`\��?���R��s]���NpQ�c1ò���UԹ�3Rx��-~�Ix��!��T��g�ș㰭�g��R{ˀ�s� ��d��l*i�Y�"�*�m�B�=B1�y�v�n4���]� f+����·9 ��L�!���%����,��@���]�=y��E�D�'�9�)�9"��LPP@���1��4�������07iȫ�f�fIe�%'��j���W�����Q��4c~`����s/a���A������I�h�@B���$G2h���q�Z<q�J#4F[g=���dc�`P0Gi\`Bd��ԛ�vĆI.�D`��p�H�c�֮\�v��Y3�h�G������"Q�^��A�c��9��L���b(�ޕ�\9�_�O�x0�?Z!�
�7	��OVp�s��=?-邼�)�|�|�ɧ�6��p��P�<w/�J����>7��A�����Ͱc`�&��ZS�[cg=�� x�@2����*F�(ܐ�.`[�zȭD��H7��k�	�HP�7a$�-��
ր{�@��u�\�
$��ܧ�����Tv"WCGX^�)��I���s��F���<��a�����⮿^���,�M3�h)�a�a���8��R ��-�VD���6��M=˛q��D(���at��(>��/����vs�k�^lȵV������]t����Xh��M�l�N�R��s���5)�u5�b�fk��'^x7�Y�{���-�1t�
�h��0����E	�X�L]v���@���Z��#y�]wu
w��\{Gw�'�~�k ��"��1*���.�p���M�A����0k�| 1���9mJ�Q���v=�G��@.Qlb9�_�}G7⫘�\{��|k�̽*Y���Z䱞C�&K)�(�<9�T����YÍX�|Q��(֜.s��	Z1TY뚊���9�Gccb����n)Sf>C`̬zy�W��o�	h��,�.v=Lk���L�؈{���j�������I��<�JY�5#��)ä����$�,�r͎�����n��ko�ڮ�/%�3��6@��G^���.���$�����	|}ɸ�{1�����<]hV?9�~_S�nLZ����g'��#}�JQ4?��.�@�e�2K��_���b	A�G�;e�κ:�Fv_W����Q ;�@*�����X�������v+&�oF�q��Ϯ�Yƣ:��g�!�cf��+q�[�\�D%�/��o�9��N�N��+AB3���G�ڳ��T%�ֻ����/7�F���W��E@o �'�,����@-Q�ܨn�1B7�-_k:����X�!@,��*.t���oPn�4�_��8C��U�PMWk�4�~���w�^ƩB��� �f���ւ��,huVl���Ϝ�'���v���3��_��v�%�;Դl�Y�{~�a�h�~�A� ����՛4�V�Q��!u���B��xJ%B�~{��8N]��]�D[�~��9��o,�ΒX�J�<�*�z^ �j���PF�1����z�Z����$]j=>�܂
��})�ܰ��G��fk�Y�%�~Z`��x�!�.����ޭ٪�ƎG���(b�F"y�ǡ�jA�;��?ޏU;v\ ��j���T���a�P�T�-�|j$�
��-$�����I=�V�dyޠb�8?GsI�~xd��6��;�`�dss&�Cjj����q6��0��Vb��n\
h���[��A�\G�ӽj����g�IQN;�(� E�vt�u�e�[	:��a1x����(g߅`,��%�U���<!8r��hR��:�"aD>lg����?'��6@uQ'�Vy/!�'��y{��n��M�=Jh<Q���^z�mǚy����!Os7��g�$�ߒ9~o�Er���=����q4�`vZ)��_eG�Yՙ������18z��i��C긙4\���9w]/G�Л�mR�����`��pyn��ɦG�@��cp�^�����h���6�4R'[���F*3H���f"��Z~?�tu�}��7nN�y_��3���C`�m�Q�*�|u�t�C`�w�B�m�xrIT���6.�?��Ϋ�p��P��v�����ލ�V,��F-�	���v��	�K�� �ől����0 ����2�q2�=s������O+��jN:3BsrA~P����^�<:�U^�,��j$��zJ�6�WҸ4�/�ˉ�+k�$��lW$6��>Χ|־�5*�Ya?��p*iP���]��muQ�?-��D���P�)�?g^����	g�0b�A5��ݨ �AWP�?��n��?�gn���zdt���l�<�z,K�	3��:-pa^�"���2��&3��r�W��३B�v�U�R��2kiz�݅Σ�;~�C;�N�k�� �YwG}`9�m��s�L���&:z^�'MS��y��q/�����U(�������r����Ҋ�*�lE�P'�Jd�'TKC�\���r��#�T�	ָ���F�����I;���3�C�ձ���v?4����/0�j��x��IϞ�gz�頚KbZ�C��]؇��!��G��d�g��[w�i�1�P4sݫl)o@�c~�^����d���H~H��
�ߺ�٧E���� w%T���7;7&YU+�n{�&y���k�J���=����.%��*�d�����۸�O�2İ�n4>n4�:Kt�/ ��[X���x*<����6�R�iQV�t"�)��j�����;��o��XsJK��Z�M#�͆��k����g7O���fkV{��h����H���0u���{�l���CI���6F��i�
!N�W�ˈ||�$$�xYV+�ȇJ��U���d]v�+Gƽ:�YM��#�#	�.���{1���@�;0X���K���0ٝf��*��wb���#�k,�����l��fy|9m�f��A��Ja"]����I���A�+4o�3U^�q��qy줥������J$SDH�K��2���w	�Ĭ�	H�,��ޫ��2�S
:�,��.{�
A;��Ea�O�%I�j֓�B�n\u'�6�u�zؙs�G,"KA7p�NMF�b�=�)��|_0��r���.e3�L[��I���_O�i�iq�ਕ!H�uXo����?�	��B.��@�5��Hg,��o�l_�d�ы��-� ?%���
'��>�
x~��5SZ��1K6�������n(���1�a	^�x�;n�=�/�Y�C��<^뵆-��g�Iq$O�.�H'�f<��T�Iy�r�޺ʝ�&���~ U�?��K2ȴ�k���ٍ�S�.���r�.��7n�R�]�ݰ ���������b4��r˝� f�k_�@�bt ˉ泒�5�(<�u��'H _9�tc���s���&��x�U�KBHL�� �y󑤼�to��I��l����T����b;�G Jn'���a�n5 ��,G� M6��E���|d�������1�?���Z�T.�Q��N���Е��>��A|�f��6�� ���،���o�U\��r�wI���K���q��m��0H��?���![c<=���%��m~�kQ�7M���1o�����e�XQ�4���Jm�_�������l4�*�$��n$��0}xR�e[Vkq5�H��������ܡ�aeMO���M�4m�|E�
]r<�A��A��Ƣ����x�l��<s���� v/X	7��:�#f��M�8j>q
��nx�FtɉC�#N�bR< �4,.��u�x���:P�vqQ�)���V�����6�+�����Aҽ0
�� �-����p<b[�3����<"G�$��9.�#:�T 7������s'�3�G��e_��)�/갼��.�<薝5(�UcL�BIe	5�$�H�EU�z�\� �)������6���56�~�s��:�.
V���ǒ.�}���V޳h>^���ɼts��e�f�c%U<�32
�͜>q�!́9=
�m��!��U$e���Yu�9X�z0�����:���P�L,QtL;��BH���U]V�ކe�=�㦛�K���N2{�&p|
@��lH�jZ����(�i�Z��U����:B�^i,?ߗ�V&�lPxZOH��::i*~�qM.�'�N���D��9�^ߧ��p�8�������]Ɖ��R������� �)�>���v�|�Ø�B7 �5'�'������'�ԍcW���7R�|g/�c���߬&0����d@T�A�O��c��UXў��J��ypkm�p9�2!D��~I�W�w(��T��^���Y{t����!CH�`[������h��V�\J.�@�)!�1H��o2z~�f�3����LSp���A���a�}љ��pp�>�[�K::��l��mj��\�L���W�N�U�{Je ���B�8>U���eÈ_��./e��`5v�ͳ2��h����~���+���gi�a��ϳp�*��N5$�[�U��(r"�C����Li��B�z-	��X�w��pc��Ou`G�i�qW�N�qXR丬�$ r�-���<���{����^-~$�`	����j��~�z`׫���eJhJT�#W�9M��[��Ǣ��,�Fe#�̵�'0�P�S� ��Iy;�,Ef�~re�l�^�gا;���K���q�A��[@Io�����{���#isT�[�|�;PB���V7ވ7|}�/])HRH�E�~6��8V�w��E�l T��Y����(b��.�ܱ�V�=���cPr>[̜&&���'�v:b�D� |g���}}�:��N<f�8����ظ��Z��T��Jɜ�`�xo�Z��1��）�n���{�o�lE$9vhW��u!vf��A ��Jy�������4����]W�Q߆�G��4�A����C����,�S^doty�3���IN0�`q��]�Ɓ�ͅ!�#Cp�z�i!���<�M�Ε���}���?�1����J�����K�\�v��py�u��PN	�
���̎��ou���*�8�z+F�j�Z����0@���1 �H8��9����#q!��&o�2ͣ����#1��K��u1�?նN�z��X�渞�w/���'kLK��s@� Mt��apgE���T��}����Um8�]H5�,��τfp����/{�����_�N��2B��#��9����V6�����)�_w�W��BGa�H�mIh{���UPC@����4�F�m���<B�>!�K��H�h�����]��6�ŏ���	��cD�h8�Y-gG��HxPN��3�>���9z�� f��A��X���o�����Nu;�W��OUΖ�[��ahヺ� ؎��|�f5���e���m�f�S�+�+�[����` �s[IU�ؼ��Y�ѿ(�M�i���:�JQ�$v�=Ð��kV^M����3_��ĈG�:.�̽��,b"�6*�ʯ�f��5��p�u{.���<�_@9�E��-k8�Zߖ�ɏ;J�.��T)Q�E���k���#._H/8���794��-�!��=N	� ���N������GO
(֍:��'�1����*z��y3ڽ�H�:�_�쬽HG�VN�xK N�е�-��Rx\[�w$��tg�������k7"�E�h5e�G���,+�*��F�]op���50��b��-o/�
��0��<1M�G��b� �&��ua�x�T��+��&9s� �#� �_R��@:�t7�;�%P�Ҹ.L��{?#���+��#���^j�e�#U��׿�9�/ȸ.�=d�SD6��S`[Y}���vq/���V1�:���r٠�Z�׉��;/�eD���cb&�4�qo��w�G�j���N5ʧR�b���{�2<�ǹq:B� o#%ѯҶ��{��-1� k:-ܑ�fiw �^K̙3���`N���g�2Y�)�Y� ��N/R<�خ�y�%R����όt�@��op�#cȄ4�N���g�{�_9Y�� [V��fĶv+�����ֿ�3��[�3���\����ݜ��
����;Y��J��Zk9���{����>T"�;#o�PfS�� �u�#�RPW�g�s̹8��)\3rΧ�(�ウ�Pւ�>l(b�[���/��k)'��W�MDOm��'zs�&���n��� �r��c[J,����0^�J����R�(x�d�Ԧy���1aWݴ�j��$)K΢8��x�>�����m��T�t;w���^�Z&�y��YM����T-�_�����L+����As��S��Ә�2x����A��Tl`ˌ�Sz�KT}p��%�N'��k���m�z��eg!&��|Y�����ᴚF| �j�$fP""z���?�٫�<H���+]��瘙���ɴť��ӯA��=�RL_�����?�=h/ds	�&�����{9���[�S�KT����ӄֿ�F��U���e�\#��/�i��~�BS��E�9�f����������kC�܄_���7~5%»�����Ye���B��ÕU!�����Hm��`:h�ė|��P�ֳ���E��3��ߧ|eUU����<ف��=,ڗ�\j���4�X��d�qMi�o��Nݛ��{6��X�׵N�(�,��R�k�z}�ɧ]�M���]hӐM?H�Sj
��ԕ����<�D�)(h'n2��+��k(�uN�w��2�t���\���*�toVړT˾�q�,FM5Y�Zh��P��W��z�<cw;ߖش�
���۾�� ��������3�L�a����ڼ�į��V��eՂ�����RM"D��ka�G�Ru��`�~̤r���֖�rQ��[�?�QƧ$E�f���_IJ�Y�����>����r�LM�c���� :E5ې�հ[��ݞ��V0�o���Fe��-,=������'���p����q��E�r���"�+��la�7 ��7d�{�=�ؐ>�,CDbW�P*m ���T��'��ݾ�h�u}K�H24��BI/�O?L�J��F���R*܃>;�dG�Zj��f�>�`Xs���1v��F�2h�Q�Ǆ�U��`�w���J\�^o�t��Ld-{2X+,#��F� �yt9 9|���h���hz�c�Z��sV05:w�Y�T��`Q�w3��%��=��X��P� a_�*�]�+�c���n��P��G���'=~X�/v�P��l>̄�>�>1?g��'-�cLʒ~�!��.,X�0��Z����YM.�
���-�@���}�n>mB�-s��~���&��`���Z
�#M� �WU�*��ꙹ�ݍ���f���L��V��W�jHj2��;W�?N	�ž���υ��j�<���V���"'�9`�  �������(�Lj.i�A���3}���^�P��r�����a�s�^�c@�ޞ��'�Ig�����H�ěZSZL)��(����A����� ���8���ri�%&	3@Ѝ2���J~�8f��e0��}�[F��s���`y�蘪�����&~��^����o�+��T�����l։�\�����W��̂���%OJTM2RB{�n��(����Wů᎙����P��	C�c*��;��m����4uH�ģ�a�Ӧ?�b{uD��|1����joL#-h}'�R<$��u?��*bqW�5��!�� �(����t񎶓Ϟ<Ə^ˤ��ԥ1��k;�?�a��q #y2!XR !0���e.7f]rM�<JP>(ˆzC
��p<!wI�{6�
I���Uߊ�r�s����Ը�u:C���h�����mT���5�\�<����D0�M�	19͜��F �����!_`OS��߿�(�l���4����}�Rya�����κ.g���Oy%�N�7���p�6�p�N��׎T{�w�.��+��t����&�@��v P�X�A}����7�d�l^-v�1�$rEF6���P�~��g��jN�(�
[ũR0�XXc�F�^�2n=�����#5��~
�S�P�vQ����׃�\GaY�Jv.�_�yX�w>�`�ݡ���؞wh�j�n�9�!��ɛ�,69���/8HV�,Q�'&0��q"k	��ɴF���+������;���D>�O��r�y~LU���؇C-f3�߾4M�U4�TfZ�?2ÝQJ`R���L��`"o����!ь�B�I�?����&��hkz��6�J�W�-6��+?��=�jaW�um�i�d�[Y�%h��
)'pC��ļ�>���QVͶ?z�)�'���`�r���jk������(!���C3[�.5�QA'��V:ͷ��R%C:4�*r���Z�W��MS5/�f9(ܵ�����+1���,�Ŷ�h�-9��×�WY-@_^<�w�2�Ž�#<
�g�$X=gD�}{�V���;�)`�b�!���n&�
�靅�?��QZ%�r^�NjӴ]N^�:X�&�M��2;+�s�Uh����,�Ü���G#���w�\+���t-#��Sض}B�8��q���DMlsW��Po��x���J#]����Q��bMՑ��D���}�)����Yp-�S
�'��U�D��72�0��K}�r �$ڃ�xKJ[8��tL_��<���x1�9*�s�/�o��z~�Tw�^�g��Aň�ڍ�9�h�4m����Hہ�y���+�����yǐE�9�B,RXPme�I+"��V�+�Qt������Ul�kh���Bpɤ��g{I�G�9�Gg��b-�,ҙpv��ҭ���r�)��
=�C�BB42MQ�T2�YS:hy|�~�.,��=o �K��+������r�u�N�rs�F7��N%י�������d�)��U����8�`Lȭye&/bU�h�jZ��]��dޞ�)��#�._1D�0Q��ޭ�c:�jY�P��J�4X�ո�~�!���TD����Q�%_
�1�����`o^;�5��%�f�]��Ž��/k��uW�&".`�*�#�Ю�U!:>���}��owG��e��$w&P�5�Bڙ��A���6�[�e�ܑ=�+o�h����jO���1�T��k��U~,�K��4z3j��7x�r�ŋ�ߏH�Z���9��������-�&d�EcU\�+���֢a��:�_� Y�M��D\/]r�?c<V4���|��o
�4c��I"97$���g���uc�=h-�e.̑�� ۽�.�>e���l�p\8pޙ��u�+�+
��/MP�wk̂��z��B��F<�ݤ*�D}��-$�_1\ee�A��q�D�����Y�N�J{%�B����aN<&:��^uŌ�-��D1��Q��� ���%�@G�qAZ�k�A�c��+�i&"�yq��U
�-c���sِ�Ãu�0��-藨�%�帝J�v��[���\�d(ȅ����iфI��[�jJ{�t�2��D�R �Q��H��@U#瓀/���1H!��Ό�^n��K�v�h��Y+��� yo�A1���&�<Nu9�}7a�t8�g�P�p\��5U)cUD�T��)Ƿb2���
U�jnw|짅^�j���[-�()�)�4&�M�[7�r�zOB�Jcd��ʑ�� �7,��5ޏ��[G�9�B���͊^�]I.����{�%��,��VݱQ�"s�������Y��	U�qy�>�y�=��oSS����{�@�)�E�9�w{?��u`@���@+'�uiv̈y�R���s)�H0W��M�+!R��D�,ί6J��}��$_�=i��� ��^���j���j�����y�

ӕ��~�kx�K��`R/yf��U;Zʾo@����8����M���H�Q����}���숦�c��;h׶R0N'��^ז7��ρ�9D�F��2��8g-���8_>G[��"r�mX;��qQ�bTlzi�^�MY\ދ�%��[��)�^�������b����ҷ9D�s��v�B���z�n�Pe�� ��9ˡ�'ހ�xe7U�����6����t��ǖ)�O㉲��6�y��B��G�Xk6�K�E��;�۔W�7S�f�A�]�T��@�GE��	4����F�|c�r�lQD���[x�#QK���o��=�����ߺ�dף��`�/�q��7��5������e�2��߅'vB��!Ȗ!ݪ���F�!�1b5��آ\C�ĩ�;�O����B��E���F.Z�:��.C>A/�����M����o^��W鶘��$H� nT�����\�.�Op�|��Ÿ0&.Q����4��29\1}!;�m]ZZ��n��!��޳@K���\rA�������bY�ۅs-�K��9^+Б��ծ���Q������\]�r�4�����oY�Ԅ��!�@� "(�IN��pO��)�fP�T��t1S	^G9ť-A���$V��GJ���yŗ�/+�[c��R�(	����K�*�_���h�'�b��X5}��6�j0<&�Q�q�q3�Ga��k�!Oo�C�Y��MD�Iq�TT�5��S��<,}+.�}4��Xl���幯���w'^��$���+��r�B�S«���t*o���qj�a��{�
�	��a~.��X@�(��8u���1��C�H��y�Vy
2�/F��_�������0�
��� R�m��+�����)a�ޕ�O�;���A1�L3�a�~��;rPc�V1��Px��R��ƞ��&8�C)��D��-�H�赶��bU��~<y.������㻍4˾n4��7��$���VU�oq	�����Љֶ�'z�R�&���`&\���<U�~A2NM둋o|�^�vr&s�R����L��}������`+��J�+����	x��uϏ�ͦWY �0�v�#���ro�4�_O�ƶ�0� �' ]��[q�=Q1mt� UAON墑|�Ϟ�W9��_u�S���eU�rK�N���\���[;}�����=j�*���=��<>����V�}@n�1�
�g]��
!m����q�PG��M�^��p,g,�DgeO��.4��p��v�/��>El�V\��"*���u0��R�/r���]�ۧ�xN�%\q�L��M�8�e�Ysj��T�j�y��^���|f/��}�Ee������I蠆��f�(���rY��t������3�Ő�7�r�$f�F������s����"��Z�4�B�ڵ���L��c��7�����˲���o�t�?��B�W&o�zJ���<�gn���ܕ2i��� @�����$�h�Э"�Q��~��%ô�XV� X��KqrI��g�!���2�+�Te9�L��߯����ۚ'9�V֍���zH�/ �+i�k%�˯i��S��ׂ��'�I�}��߆�����[�#��yu�����@�ǎK���٨+̓?ݹ�ir���wf�D,�8���Q(��Oea��.�ɯW��Xs��Gd�@'�d�Fb$�苎�>a.R��������5$�&�2y�m�^�
$G��]O�Ϣ���R���@v��jz��ٓ�f�1)�FiN?�pC|��Y�[�O��sS��� ��O������^-טs���A�\7���
���]`�����l��5�Q�n�m��-��0]ݣ���ˤ�
m��E��;�ѐ�ץU�C�V��/�A¶�%��L,O�ȭ6��Q��3�<)G����W�4r��h��OzQ�a<W͟C2*e�I'⽥" �Y���&'ĿeW�;,�k�ų�8��ڴ��.����΀ffѶ�-��B���C:�Ti�����ȸ�z)����N��7�i[�Ґ�J���Fd&V�u� e����- �k���M��VwD��G��l��M���q॑R����I99r)���f��Xv�F�jX#@���7�
d2D���1��q_�ʈ|�,�d)��^�إ�aY�_��U�ZhHP/���d�&6�N��ml���m8�P�wa�0Y5Y�v	+�����E��W��b[���[��q�B#D�A/�j�0EO="�<��T1�iV��S��] P�oh~W@����;d���ʍ�bBX�[�9�+D&���x9<��s@�{��B�K����QUQ�k7�s��v����
�G�?��G��+��
�����&��������G@ARv��k�}��>���a���i~m���z0�Ԫg�㍇iL�"xm	N�2��<��aI{M�-9������7���^zRwΛ�q;��xd{a�9���ծЅ���Y>���õQ��7�+6ɔ��V�U������2�\b���@@	E�8�O:_�e�xvp��&�\��fW��d���/�~L	�%����3��J�&N��iʧ�	�"�=���΋[�tll�G��6c-����?�=DF:��Q�� x_	#`�P��3�9��GEI!	�/��GH5�X�l[^@\f~�l����tIq���DR��m9@c`V�8&il��2��Z"��髦���?�=rTK����0�C�H��908(��p��a�`�Y>6�KZ� �&���ʣ��F�Y��5x��Y}��4{�ĥ�A�\�H6�#^s�Փ�>�;�˕ � ���W�|-��x��i W&γ'%�A�n��4�� s�<*��+��)��wq�K��
 �/0<�JϽ�ڼDsQyo��1r�S�j߈�\k���rwx������U3u�b��wU�r�4�oSQ�c��=ت:�y�!*A̩R��+t�Z0_ł��3��)hIN�ʅ:a��=|��CI?�A㆖�����Y�c^�e��ƣ-ؓ97wB���T���^%Z.�$�H�m�ע����XF(]�VP|�W5<�7���/_zk$��~<w����4X��"��B�ث��&��(���*JF-3D�T`6L���W���2�������]4o~ĨƂBc�,=/h��~ѱ�����5�AY0o����b��wS�h]�'�O6��4K�X�Bv�
��Ȁ�x��#��̧j�7u����1G��iB�@�F� ����-� ����F�&p^����-�2CG����4�V	�
���%2!��5�غ[3[����9�7gA����T!eS�x`T�A4�=R�]�8�f��I�O�4Uءͣ�Ԅ<0�[�ƣx4��*���3����(��Z�p���� �&��営J�H+�HɟL��D�T��Y�֝�t�٤���o�Ў��'�A^M걏��RTǺ��|���R���[�|-��cu��p���6<N;'zP����lv��߁�3F���8L8D��F
�_>�ܐ�c�:���ᎈ�Dh���j)+���d�*W�����p��?BY/�)����������@�mx#c���l-B�a8"\b2�� W.�9������詧gVŞt�H�\~�°z���Є�fׂ���98�W� �z�N�W�S �|��ޡ�
"9u"_Y-�c�:v=v��X,����Gmy
;i3��_&���AB��Dz��xQ	�`�y2@����tp8;�&�T���Y~à� ��hфq��gE�L��֍.�W��25��,�GoV�o[V�7�n�ձP)3s,�ޡ���Uzt���7��P�P����PEf�.�4�s!�j�݊c��B��f0B	�бUO��Le���L_��b���5�Ϩq���P���$����\�v�.Yu����H;��C�>?5�<u�q�&��Q������l,=�[���'':WS�*M�^������������+�pQ���Q#���^�G��K׊����Z��z���:z@����\d���x�<��}�k̵W�}��${-(9��o޴�ѱM�()F�Y��ê��$]���Z�f�3�#`��O�:�;�ۙoq`�:=EiG(hU�n~���H5���ʭXj�� 1^y#ݴ(��v�*�x����XS��{Ux!^l>��'���d�W��:=���p��\6���\+�F� i;���;5��ԋ�^[��A%&�_�+o05���z�Z�µ���|�YH� ��${��ä�2�d ���L4Jj���<�wa9ѫ���*������5��٤%B܃Ǽ:1�:�����汲�.�W6X��X�m��8{�����cF|�NVbt
F��8�D�����V���A��\�_�6���|���3��3ô���^8>E�����I�r}|F�5gC�I������U���C;�%Q�S���ȼ������O�b���2�a3� u�k�_!$��ݼ����>�������������O-��J��
��;��Wb�pe�A /��fRե�+�����gZ���Џ[|���n�AVC�B
5tc�ɪگL�U��Z67}:V#����u�qS�-z���2��NÜI��m�N-�+˿����1I����rUoU�7?R��-�ګ�������Nԯ" Ћ!��8�c������ [��qL|��
DU�m�O��A�<I��#3�c��s���
+"�쬎F�=�x��5p�(o���� *� D7;CJV$��[Mm]����.�e���H ����nZ�*X����??*��ޥ�NS�ڸ��?��_DƯp��G�t rLl�,j,T�J��yj?�8B
����>�o�W��ޑ��J�L9�S~RW�.Ll|"z�?�$�ޕ^���z�S*{L~qe��xIJ^h&��2�ǔ��L�����n`pQO�վ�j㇇���� Rs��ߣ�an���4�A�k�jU��Z��<p䈳����R%�s�w�@�Z#���	�{��j~G��0CQ<9��˴�]d�	�W��NY�Ss`��-Hg�:%��n��"��8H"g%�7��#�R��I;,�6;&�
������L�"��7觡W���ӛ��Y"����yml�i8X�
T ��ɬc��������{h�ݗ�u�d��g�\�)�~�V�X;����_��Zw�珞�$|����2W6���`65�g���FM����������I�ftFic!�Fqn���q���T��r,�$4b ���n0�? qɮZ.����`��`d���7$�0�m������I��Q��>��a_��9�j�/8�a����\Q�7B�\�(���D�Q�_�/�Q����d8��6J`9Ĩ1�1��<��+$��xbN㑟�h��]�䵄��|���)���Lf�v| e�Qx �19n�?Ӽ�x��A�u��6y�.:N6]̖�Υ��^�� �f�rPc���X��u��#@&c_�s�m��s�Z�3��6����"�W��l�*����嵀���5���`����Eus�F�A�I`$�F~A�����Zﴡ�Q㉝���=���`��dU�H��:O�0�6[�E?�ւoo�6<PS�|�h���,��E��D (M-�)��U�A�Q��4����c���.�_�.��\m�>������9�J;����M���<q�7p�����#9�zQb��P	�h+h��w����uׁ���ˈ���٣=���X��t�b���E�o���;�qaoƎ~��f�,i��1�.�X�T�L+���)��)G3�A�D7������S��Cŝq�2Ƚ ��6.�v�+�"������A����^x�.�fAr�}U���{�(p4�Cʐ� ���FZ�U`�������a_����n$C� �('��C_ٝÞ�h�׳���<���,|��"�����$� Wj�g�^t*=����u`$C��0Q��t�Dp���p|-�畆��ϻ?���=Q4{Ԙ»����D�(�Ǔ�[mV�l�<�Q�4��I�B:�E�^~O�ߩ�k�Į�gJr�$h���Yҹ��B�Ad��"���f������2a��c�sx��yKa
�v�NŃ��!��v��&>_2�tZͷ�i-Jt�VL 9�Aไ��y��H1w��`�Z�<�|Vr!0}{�u�^ѐ��\�$4:�Jd����`Z���S�mK�� ��_�/��M�|z�g��s�$�HҪ.j��	�� D2�ǾU���@,�߳�ؕ��m��8$a��M�@50T�-&�'�{�w�����ZXKV�����H~��@�[��ה�W�{�}��]��p�1�\z�eXB�����\+��]�$�
n�1=-a�W1��@|�������MG�����e�;�9����Q^�&n����l�*�08?���*�B�:������fOƘ�V�c�-PY�~C,��Q�}���� [s l����K����؝�qc.1���M��c�^�`V��uI��u��/5z"}��OН�`M�.�t���ui�v�&�H��;�6wC*2����z���
����9U����a��6EW����6+3I*��~�t���4jP��s��J٦��۾�[/mN�N.�nX���WuN�=�2kY'�-�,��q���^ꁲi��/�E�yR��gb��[�}n�P��tؕ���D�X#$6NGR叀��t:����\�M�B4N���wc+�T,��|���zkM����MV�پ�sA6��Mz|�T�7@ٺH�Q���b�}W:�������cU��IjeνMK8�i�ү�A���P���h.�!l2'l��r-����4��,8�	ǻC ��h`���j�5�NE�%`ѪG�S�C!���K���[�^?m��Џ�5Ϥ8ʲ��^G~) ��Ϋ���n����ʯR���n�&a8���&�	���@���(�Jأ"�oT�6R�v���|\������6��)�Yq��Q��=���0:Z���f�׻��Y��L�I\v���]�z�{� �g�N�p!�jf�2QJ�Fx
��h��ңr��W�#|.��R3)Au��s�	$'d�|{R�iR6�����K6:.�Z��5�k�py,���"�d��Zg�s��ğ������kw��6,�����c��-_9��DT����Ӏ�oy(0>����f�E�c�>���`�@�n}`�X��j���/w,.k���vձ�WZ<�S(�[A�TWf����L�O�{��6��s!I� :������z�@L�9b� �'R�Wȁ� �}�!XW��Eq�=p���>YG�G���|Ճ�ۚ�r��������A4�V�)D�'����BC���b���h�;:#y��@`}1&M��X~8�`�e-$):����Ѭ��F��_9JC����O�/���	'붻�9�59��V�u���7K��x��v�Z�'OB�:�����_>���&�����,�{M����ވ�ÿ)s%c��k����}?:����F� ����]we���3x��G��B����4/�M�����ӿ�����Kw�}i?���m�n�)x7&V�)`�8�,�KÊ�.�XJEɡ�f�;*<��Cz�W3�g����*Ώ�,�MY��QCG�2}.����,�"͛Y��~ X,��%���)x�<�!�s��OJ�	�c7�H���x��!�pum��~%u��Wj�=Dd&�/�E�-}��C�]���evsK�D�����	�@(��D�ste>h]�����$;ܶ.Tc��E.�:ڳ�?��&_���aՌ��T����,l��*���x}�L��%���p�jX����9~P4lw��ƠR�_/�݅ �����,��cۭd���{'v/ ?/{ǋI+p�wʈI$z�QW���:/ה1�~q���%2w;po:XC�@@#wB��4��`���mh��U�C	�vp�x�Y��EC�[����$���$B�y��c�r3G��dY\S�g�Y;7���|s��q�zA!w���pKs>%�2�)ܓ߃�+.ٟ�8އxp��l�V���*/:l��e����{��)�'�;l	�Ŗ(��w+��F�'�]����}_�)˲����{Uy�;^�$�.0s��h��_P������-�>3a�Ӿ�B�>�����&0�8b���Ӵ�HݥF�Rz�L���]�r���b�Wmh�g��:.��т�vR92ӈܫQ�
^䓰w������o��-@S�W⍷_Q�����KI�|�4�q�f�����5p�x"���t���������]�@��N~�ak��Ѵ��}���4����ê�rqe�^ ߚwK�f�e����a� l<$,��)�լ�>��j��3Ӗ��3/�W�rF��:y��B�-�j���CE�c2���W�E*S(���o���Th�����aY��!En�14�p^�ץ�Tl�6@U��B�K���P(����fg��4��,�2�zf�]�l����^����tM��Ah�Y�y�����I?I0)�:ܛ��5l���u�~�e�УK��NDh<4L~�T��5iڞ�Х�w�H����(nئb9$M�.��c^֗�kdd�3����R�,?�O� x�[��N�}�"��U�XT��������C��[�W�ɿU	s�{jA�^z�_���gj��Z���O1��9�e��1e���V-��V�v��.���2<Aߥx5�*�L��5���m�Bp��;��t����47Gc��,Q�|!�m��[̮J۹C�ID�L	�nmD�NJ�R�����"S#�"FC-��h>M�G�Cڮ?W��ٱ߁A�� ,��:�-�-��L�'b�$
#C��wNy�Q�U��v&���&� �k��ms_�*
�՚�+J����y �}k=�úV >���+�:R��1
wA����,_��m�Hi'9���;�~ vO6���P$��9I�Žz��=�L����,�uQ�h��#Zf��E��i�L:H�7aD* �A�.2�#1���O����뼔��s�, /��vM�q���.1c�nU��c��Bl\�K��~�iLL���&���p�"v~�78�ƖC���vOv쎹G���;�$H��u�pM3ϑ,�#d&�u�`z��B��G����A��2���#t������=ta��R�ߎC�d��o�Z	5a���|�X�X|��3dT��gN�,��w,�Е��'U�6QqPӜ��Gv
�X�Z}��t�����C9m�{�ط���8UzbgY�	�bu� �|���hPm[���S�uN����󈑵����5�3ŷA*O����%�u����ō�R� �E:�;�܀���5��e^��a��НQS���N*� }��LKz>��s��cy�t��ûʠ޺�������S���XU���p�Uj髲�R2�vE���n���G9�K�TM��x�x��^��"�(1轃��K�+�EWm'c��b|����/��B�=���[C�_3#Χ ֞� u���#��5dg�X)��2�E���B�YZ+�%�T�>C�Դ�����qG_��b|��/垉pL�0�s��}4$
Yo�b��#�UB(��73-���p����*��������ЇS��p0�M���r3�Yuƍ�x�4�>��]H�M��M���yp2)��px�=�Q(!f��8������m���M֡�J�}�xv2Ѥ|��LW,��ǅ��3���z��ϫG3!��[㬖�O�w����Ws��H�*��E5Iri ��
OUe���
�Z�4�*����T��**M��U�q�V�M >�Hu���g�k�0�W�cQ�ؙ���3e���~�Q?��FVH�����p�����=�}ϱ/�ṍ߽��w*�'�����F&�C��Z���ђ�$h�lM+Y�Z����@��J�Q��j%��ޕO��[�W{�U/�Gw�J���${����3���pv�搽�~�J�AW��Mۭ����w�Y�ieD�֎*6ܨP��_r �h;�X����X�<��`�ϋ��9꫼9��l9��tGPİ�ӥs�2����ڽ%$�V"���*ߍT�7ڷ�%��-�g�蚡��E�-�b�4�]��-FMOz�+�O��1C����+�����0�̃�.k����C8s�!�W�� �H9Z/��)e���T����r��hu��0�h�;E,�D?>���f��`�jůeg�Z�Z����4�Ԩ(�v
�X��u�}>�(F�� 	�וܴ�R�`:�� ݀��k,������8��\��x���M����A��Boo��?;�K���̖��\�7�7�@�-'�˫i݄w�0�A���'�'��|�~	+���9Ĉ���*���T1����פm����(��Q�% L�z
e�<z�B]X&��a�vʞ�=n1ZE�U�,��!�R����~��R�����V��bJ$�.f&6��4`]��APT��q��=����P��P�h�T������)ц#A��1���-�%	���cd}�}���˹55��3Gܐ���A��%�^�8xBl�7���q������<�����A�~�~:3���4Q�-���Ϻ0��r�jn�A!z�6�?��J��[�m���>4����O?l9c[�"��f?����5����wW�cf�6��|&�Od�}t<.yL����1f���d�`q�vH�хt�oSW-c���?�~�-?0e�x�_'�U���M�	��NmGDl`�?���/S��_�2F*�L��J��V���сi?�����԰��v�bu�h�N1Y��8�ϯo��0u��d������B��M�w��  �-d���^�wj"��K�+��]y�^,�HȢ�X�@i�{�I3x�a����e�L����������T`��<+������EO��ӯy���.Ś?q��c��]��v�\&�ԧ�X�?��s�a��Jj�X�h&<�T�I�n�@J�EN�^+Ν���{���s����Ԟ�X	�6�obP݅��։x�w,�f�����R݃��=�(���Wկ�ϴ����Gy�`!�*�I�	�(�r�P`��K��g+�H1�䩖z��J��/§]�eu�v!r'*�7Ą�~�4��F�0`F-V�O7��r����H|A#����H3��: �~L�@�����|ହ��̦A�ĮO�PPvi���Wy��#J�(�8�W�u�Ǵa'���Qnz��ؔQ;Љ@z�T��)7���$d� ��3�:�n���P�6Է�k�W����w0^�e���oWݗ3%q��LRh�x�&��yn��,�(w.		\C�S���gw:����y��^�
iq�Ҙ,����&��خ�����C��e�m�g�ͩ�<�C�B��
J �e�_`81��z��HPePP<�j�����S��{���w4O۶J�>���헾mt��8�I�{��ߦr���Cq�_�(%�� ��\�H��u�4�jW�
��	XI=�I���O~ Z��w����+wSg��(Jmze���xY�8ջ�.�`�Va{��L��Y�]
l����滪z�������ʇ�1�=hU���qX	2-���]�Qj3^�:���5m�P�9B(��ιg��n�0k�rL'Qv���%���H�Թ�ܼR��$���$0�_5
����͠-������`� ��&��Hib	pۣ۫Q{���e�y��v q�N&tD<f��_��1<�-�ga�z��;�.�E���r���T�OH]jZ�9��lO��;�þ��t�Tyz�m�1��_#ɉ������_�A��:���\�K��ĳ�->	a���t����F:��}U#Q�i#��KS�^��]�n�Qy���U]_L]]Uߨ"K(ܼ�$�,�s6 �����\��f&�3��!�J���y���<ǱJ�.�~�����F1�K]Iq˰�kn	Fw�yd~�-�K�Q�8�v�4�a�.Nҋ�U�4�Ѭi�}��Ũ�/����q6�o����,�q��������$��ji3ڠ�|�LCg	�z�0��!޼2}��1w�J!5c�bo(�4��6�/����>J�x'L[�[#���΅��Xd���1�@p�aS���齶�VYlɊ��TlQ���H����!C��k!�?@��V�o��G.^Xf��U�=�gX5�3��"w�G��zW|���ɶ���M΍-�>R�h������P�ok^��d��:�����;�Ŋ�z�@6��c<Fo��*ٞ M="?��^���*bc�A��<[:��T2��ph��-�1�����!f�����R ���Ƹ9.ٝy𓜰����3#匀gv�b���l�|v&H停r��j{�f��´�
��̭4>HW�ꮛؿ�E�o�c\<�7q)�	e�eZ����9L ���	O��QL������t�5��Z�u���W���PjN�r�)xGo��'S�U�O���[�N�,��\GؒN�'*�g�Ϡe2��E�O!�����Cİwcg+�_V���^'W�����sw���4(
�)���=�t����D?+���k�LPQ-���	�=b�~�X\�J�T_���i�eZɆ�Q��ȤU��SG�~G��D!���0Z�z&�YLl[���E�Ҟ���7%��'ot�jR��k\���6�F���nJ��/���Q!@�����R@���~v�G�F���;")n�%��:�E�֌F�=a�Jk���s�!��\�nncE8�O'���o/��R��Q�ƿ��%~P���.m|�֖����tuҝ��z���kTګ<h��k��q�|��-�fW�\X�Ӧl����D_�P�D��Aw,�Lޤ�tow�*i�P�R�_Kbf�Q����F��6�`�i{��Z�+�:�I@���X'ӈ".�"IE,#\G�\��T��,��u��/���Q��
��ɤ��}���u�:��/�=X͈�������h��m͢�HsQ�Q0�H��`N��-���l�<�G}� %v�yA�n��5M����	��׵��`�z�����_�`Rs���'�taG؋ii;o��L�l���[�����w2a?䋜��������O�L��~�:�i�+��%�s�Ϋ�+Bѱ���)�V��u�[�٘�*{�40�%���U���G�nK��Ht�`��_.�1���Z��jG�G��:��?�̯���7v�"����c���F������"��}�L�ʧ1t�R��;C#7\��f����(��Q0�ې;��S��� g��y��*C ����|?�m,c^"���#h"<�V�N�k����2^IkT����b��b�lF��&�V
y�d�8���aH*W�S���X��R�@��Y�Op2���sq�F���$�-�.���E*6��`�^6�H�����2���k["k������`��}M�Oe1��IH��me@�)�>��@?�f�g1���I��E�lR U�����QT"�I��to���Wb�<bCHV`-ql�M��������tV��us
��j�H�=佐� ������ �h�������@��p��D�}���@�-ZF)}�R�Ć?V>�	��)�����{x2�"����lc����Hw�=�"��J�k�z4m�5��	I�a�&�/�;�����֕	���naw�)1��ĥd��ş�*�� E��ޤOs��a�˨9	��D��tX��z��u�|���N�� �3�%�ז�f���*�l̵��p���H�{�ou0�C�{$��G�O@�7�{�He�9� ]no/�u.�:�����L�Dw���%���z'��w�+�-���p�G�B��hg���
�$iTt�V�u��iY��W
��t�@��"����u�f�R�#��՛k�i4_�P�S��eXk�N��!�۝ A�T?�#���E���Q�_�
wL�[���i
vYk�hhZ��g���pK�=�l�$̭͖��l�V���՛h�\iz�/�pA���20����B�8N�Q�G�55�/gaF�H�2����ɪ�\'�V�!~�d.��|�˸ʅv���V����ʂۊ%	=����yr@2���Q���e\��C��($+�
{g���7�&�[L]����:M?2{jN<�n�/��������T���;Z8�n �_Q��G��L��*ʂ'�'����u]j�J���xG} 0dޜW5�D���0y���{
�B�S{��c�2�󷑎ק'���B|%�	�:dl�[8�GQ�B�����"ꂃzD�Y�e���Iw;=b��h3�O�%��.��h�qk&���5vl��V��YnA���(4�1�kyY��bd�@ ���U��Rni�(�Y"R�+*�v����ۭ��"в�*��ZM�e�F�h{�]��[{.갆y�T�=LL��c\��1�Z�/�>��⡧����#�+�K'�"M��nvLҘ%Q�e`>p��dW$�t�ܠd��/���F.��z��b8��L�=.�u�@cXS��Cs�~�0��
��}v:t(�n�#�����y�� +�(�^	[�#� �y8��
i�C2�sa6j�O�խr�*��%���xcx��9x ����%�|�7�d}�]��S]��LP^�G5��0q��i�����S��v�J�������[��Y�#�LSO=��d�H��*ޤ/�	:��<ѻ��Ñ�<V��t\'�<#Tѓ��ĺ5"�&���H�i<�p������z�+�Ww�	q{�^��G-��f0!�����Ⱦ�f�0|��Ö��@���lc�
uy �y6Rl��9~+SlG9�K'n����:p:��%(q���)��{�bR	c���~�����U�6@)Èo�"����(��C^�!��R�X��N߼])%~��V&ls��s�K�撲��I�t\��H�� �e"��.�)��
$'��g��jL�����֩j���G�~�j���O�;^ĝdd��%sDY�s�K\���\*%��:��a�_(������)[q����? C���Ϙ ����3�L}Ni�w����7�)
��̧IQL�J���a��.�&#EHQ���u[O��K�w���Ӌ���X����ʜ����2��$�F6M,�m_�ڗ~�a6\�N�3��Y
bhS��3C����<��:���&�.FU�������,�Ȟ"�x/���a��,8�=35���K���^*�V��r�.��&����>�Ae��? �q�����#a����J�E%��ؾ��N�ÿx�N5��jX�� ��iy�����������zq
�~&��$�� 98H�|A��Gfܴ�?���[�Hp������U����H�\#O�̌:ᚨ!�#
G����~�w�a��^K�מF��3�7.�Bm�\QA*z� 4fzG�������9\��6��Kb���HY%���b�E�wsC�ߕ�w�8m�_B���հƿ��&�Q*Q�	�x6v=�p}7�@�b��mK!�$)mf�qk�
C(����b���K9N�������[���@��=nq��T�t	�}=<q�B���\�����y}���[:����s)�W�!��R�����A���}c��HM�M.���٩����H3��;���T3��𶅹��)yW_��q'�:�J}^��R�I���[�Jx.\y�5Đ���y�p��8)Q���l�ܷ�ٕ�v�������InP�h�aKL�hO�?J��;ٱ��1=�{F>�(�ͦ�K�8u�u������߀kKX/�u�ͰB|���{�w��Q}�8]A��"��v��M ��L���ܦO��9{Z��*�^q�!-�i@h� L�0x��C�Y�&F�-�g��>>9-;�yM\\��Į ���!�6F�
�1.���~�C�w�L
�3*��M`ͣ
IY�B��%�Ǹ�k?n�sE1/�¨��~�c~�%>�p,#�ң��´��ˉ�/���J}�8��'�눏�I�'�BuqxU��ە��D�U	�=]!@�>��st�d{oY�X�YoX�b,g���P'��_�E��Q-��z�ƅ�Vo
�Ŗ5^[�����B�#�݄O��x�9[R��-P�����C������@m�͏=.�����.j1�X�:�>rD��L��.a��=,k��M1�h)�kZ�,�_#Y0S��Y+L�M/�FR�C��JUz΃��qYw�eVuR������ӹ�E�	5J�c�0^�9ק>����0J_E�g�9_ԉ�L^gW�W��r�|(�`��?�|���]2��Mz��k8ɫ�������%\ͬ���ip%bM�'�C`H�3�`�>����%�� 7�`�8�C���I1_�omΧ0�*��6��&�h���gB?��>�'�����n;�^]�'z%����=U�|��m�����W��W�=�~w�+:�]}�ȫG_�\�V����y �g���w"���@_�k>�cbm!�v8L�,�go����G��G�B���J$y>���gXN w�L��L߹�#*jifT�K����!�ا`W�'���P*���d��(����ʱ�n{V�����̌/ln1�Z0�j�G��\�<���9��NP%���Tr�"�����҈�rPi�@ݹ����_,#�B ���/�1�m����1"4Ɨ&�h�+�$/�4Z�?�u7����Ƥ?��$?��&�^wົs}1��l�H�Lęx�)3�--��cՃ��cW�B<v�܌�)�/.�NE	�9����=Os��Q����b�Fb���9�rf�DID7+w�|��V��cwvV;�.�09c���@l"�]A@	�Z����߂?��v�C�E�b���[�+C���.W2�P�a��!H9��������"#��z�$>�}j�;tP;����B%{�X"XLu0h*L!��@�J���������,�[\r;���^]KE�|�O��!�v`sw
#�2�`~�ݲҪ3�Cu-#���TW6��a&}�+��b�$�ٟW�ܕ�g�I�0|E��'���N�X�
�H�A�l���ͤ���q���$,����9�?�Q9{���p�ЃB�3.�zp�kS�x�������OR:�d���<���УjUxv�d���ǈ�+��<Nψ�U�\SH�{�mQ��D6�U½����^��ռ�1a ����\��
q�S�-��x�'F�k$�G�M+�� ��;�봮���7N����Oۣ�}~���I粦G昡��ܽo����񦡩y��Jl|�!,~���.�z>�:���r�#:�[���D�d �L��[�9A��CƟ�sQ3we��K	3䰝s�8X��0a����Z6b0��R��IZ�ԎN>N��.��Ga���N�����3Z�kK0�v��}!���-V|�!�V�ޔa��'��s E�l,6�p��[ݭw����Go�@/"�Ct ��4����E+�&�k�,!l��ȲO�V}��^�t��J7��GVjHy�*��V|n]��4p�P�x�h�+f9�5ٱ�S[ZI�#���Gs��@�QC������Y.���!�
?�c�W�:�?q�r��0r&����#v
���LP^ع* gj$��p��y9���zkd�����������e3�vI_��nط���F���D~F�7����|3���u��1-�=G�������{R�	m�U�����=��-��@&�K�E/a^P$ ��0'D��`��"����3
�L�(���@��GI�*[�/���J��p@��JKfn���Ϗx,��Q@��4H��?U�{��2�̌I�S9�ٽ#1��aĈ$lT�}f���J���ȷm�+�C�AjH4k�^}z��;�8bFw�b�&˨����0-;h����9KO	 N�C�cʁ�Fi��*���4z�&�Q(��;�g2�����*�/���zX��ԄJ����<HP%��ez׆U�8��� =�i���a�[l�j�J�<΢�#(o[�/�wlc�\,��'hޡ>a�'���|B��-���I�Sz�G�g3�ۃ,��?w�Tc��peI1LH2(�)`콋s��U��?w�h�і��&4��E��<��ݨu��0D�����k�jL���}��\/�c��2Y�*��ń.�u��ҕ�DW��|��^��B:�rQ8ۡ�^��׽�/ݫ�4�9`��f�(��P<�|�4��_0��}�U.����03F���݂�@�
 _�j<d�P���T�n���@��~���f��,��$!
mO�r2��}]���!3�G
zL9�	�l9��46R�TIq|��0'��@����<u��_�	���|�;^�r4;�rK��P���ͦ��v}�i#��&����K9z�R-�ip��1L�zdҥB��9����/g՛��3���D�ԅ
kGц+�WD�Q�g�iN��1�RX~�z�NX���m�W��E��O[�T�� �Ҭ�/��鶺Zc���>��cm�[��d)	h�4]o�!�7�k�83Q���~��:�˿v�bt}������*�D��������u!
6٢E�����z ��t#ڵm=�u��]h�v�����P�T���%)�	\�r���{��e
A�>?@%����K�C]�O��,6"�"���y�ih�����'{*#��I���W�������@3�ނ�o�eaMe�O�k�c'H�L������3-^���� +1�<���n�����Z�Xw��3��' 0I�]�>7�T�1=p�fz��i(��Bhx��8�͵dq�؅O�|�pd~WE%?}��!L�w����q�A%Ҿ�i���$�H��J�	Д�	o�OQN(�3: �el��z,���Bp��IiL�5�!���?�<�(�L�e4��kJ=,����Rք%2
x6��Ƃ�	_��_4�qDj�^�׌C�4l�4U������]�]�?a�K��B��Z?�G�_�=�s�o�a�E�g ���(�����<�l
[E8��v�'�����Y�MW����0 y �Ok��IQӅ�gJPa��q&Z�)I�uI"��U��3����MfI��/7��NS|V)��M���Kh�� ]N65Z�\��4��܏�@Y���/��nY�R�J^���lw�F�D�|t7N;|U��m}L!�E���c6��
 3���6Y1�h�ڕ��LRe�^��pї=����G��oQu�/�6�O�U�QH3��x��7�
tN�	$�Tj��� G�E�OXS�&�`��yZX>ts�-�`����*�7��w�Ŝy��hk�-c&9t���l����o�K&<ɡ��hn�Q��}���V���
�0���Óuu��f��CB-���@g~������~K�?.ɶ��E�o_&_��z�!�3�A��D9b]W��$.pa�g����Q�K*�k�I�)J$A����)	�F�p]��~���������Ah��I�AcvCH�������u��6����(̎��ծ�cg>��n{�R�_:&�@�z��q�x�K�� Q���{�N��6|���l�'3��W�o�Ey�%�]>��z���)B+�^d	���$b&�|�o�Ik;D�{���e�0mׅ.���B��ѧyŸ��6
��%��402��� jM&��,�kn�#q��K�Z %)�S��I���{qd�AL�%in�>U�XR�w�G��2�<���\�V_��A~R��&�����0A���a��qY@�܄�`h�,�5
�̀�B��a�mMin�+O��EM~-BnB*i�REh]��
�
����/�,�+���ж���6�� _�P�t�����3/����� ���pp�P�O���줤��@�"����b�|�uH�#'e�:���]��E1��	*5���N����ڋT	�j�1)L'sǸ�e�e�l7B,w��e* ��(��]����㛢�?�� ���G�C�& ��h9�h�]W��Uġ��w������� �K���P�RU>}Vn]`�i��F�7�'-UT+�5u�u-AY5?��ۙ�������u/�����Lcj�ԒZ��U�'6%�2�o�z�{�	 5k����e�����/��кC@C��-N��TG[��,9�o_d�v�f�����\�Ve�&r���z��柡g�6�Y�`��a���SJ�{"j�_��ڀa�mW�<'���vz��r��mHv�O�����,��V��b�~��"k��JJ�4�y[z������u�$�/	!	@x��f�-���D_�����_���jb!.�2B��d�<����u�W�Ⱦ�/r�(�"�pI���ꡩ"�K!>��;���ӮsLk�)���m:\n{G�E$�衞P9l�g�W���1�
0�&�h ����<�ͳ�Õ�}���o�T7P�9a[\LLr����<G�)�#'�c+<��?�p'ٮ)��C��*��G�hJ~v!���*�ù2�S�(z�&ɓ�up9qO[)o����*������k�8��vɔ������Dr���7	 3u,���&�C��POJ��B�R��^!,z@�UiRw\�D.g�����'��D�����{��?�U�;,'�{��-�uV|ª��AH��U
�#�h���Ds�%�4c�U�pw1��^�� ���_vx"2��;�1��c-6�YϦuŎ̑�n3�j"��⋳m���K�J>����ldPQ�Br�c.�m����y*����hcWw�h�[�~��&�("���-aTZm�0����%F�'_�	"�����2��w՘|�ZԵ&��p���!�@�MCbAr��s�,�Wᡸ�%�+av����',��I5F��F'L:�|� 00̞��K.w�=]�aĠ���=��jC�ܙ�z
D���eKV�m �ml�nk/\_6�9'{E(�(y=�i(�7FpX~[����8�c3S/5�u�G����45ި���p���!�&Pд��]�T0~��&��l�"��(ؽ��.$���p)c�}�+R)RJ'�g�*{���L��=^)���-,���B@�{���%R��̅T�Y�xd�CA�(@��{����I��i!�̺�"fTR�ڙLB&��u�ޏ����p�?C������R`�:͵%���"(���b�ϗ�[��s��:p ����67��������d~#$�!�V��p����8�;�t�6N��%^4ZI��V�lkuf���{�`0T��Ўtd�+���큦�f�{
��4�Zg/Bĉ{���1~-&[��m�q���%����L�u��`I"&������	��{�9�r9ض�dԆ�5��U�����S@T�Z6.�Ɏf�$1�[1�%��7��k~��fM��k֊���\*�:Lg&��Q���G�6�!�_��w��W��La=W�W?äU��h�`�.�P%^}[����+���Ơe�8v�Ӟ W��@�lx�S�Ad��-�R���ɘ]�)=.��BQd �>�w�9F�M��,���Oaʦ��/�ɦ~T?��ɔR���n����xmKv�D}@��r.��#<���q����3G��hu�8�.ᚏ'��B������;�����j	�%����Y�������No�G�����I����D�o���*6�V���#-1i�aAT1��o n-�����|�_�v�)��C-���j��=��^��L׿�v�C7#` ߕ��iL8h&�u���wB��bmq.5��z��C�<}����Ƃ�&7�<  9;&s�s�3+L�#D��Ŷ|[����m${���lB��55vXZJ"d��dqz�w��f�Tf�6ʵ����Q��}������߹Z9		�> ��yj�4H�Q�aa҂�y������'�,�b��\�����>��^U(�)4��z`��ቺ���P���E�ٰO\��-s�^�����;�ݷi|ژ��+�O�	t�j�,�|6��<��6xj.I ^�\�����m�������zϢ����V��$?~����]������H� ��u�?��D�B�d�#�F���GIpKu ��jAj!�_w�&�O��quI���KN�\���DSq2�j�-�Ǚ֫q���>�H��ɜ�yw���wOW>��J������	7ֲ�K/� �qKt��/���P�Uɸr.��=�e�-t(>���+p'�a�Ij�9�X-iM���u��A�S�p�^,jH��wG���L	��7 {'�h*i���9)kn�&�7Nۙ��G��Y� �0���n?J���lHB;��I��'t�]�3�ix�tu��.���TS��M6�e�,�[��_�w'|�y���	���������^kOغ,��d�c11]0d��|U��v�W�d���w}@�/)����a� �Z�ƉBV��x^|��L<y��4�+���2>h��/@�����x�ԁ�|��@s�
�<i�i����ϕ;����R�Z��ʔ	Ձ7�m��*rN�dJ���,�v.�VB�X�������c��L�Vu"=�������6����`TaɥA��믝h�JrN1m�Z��b���M�����R|j(��/!��ا�����)�'1�Z(�i�$03�qk�]a�.�����j��J�`:zD��VSlE�m܆D�~���5[Ej�1hӬ�2�Kc�n�҂u�i'O��00_S�����X�q�������Ls=� �#��ތ8Ɣ����b����//����1٦�{��ka�c_m�H}탦�}����h��A�Ys�Q�p	�%l�WiP���2���P������ǰ#�蜺[=���8Xf5����䨭L:bj�e�R�*͹w���fWu�m�،*OFe-�� k\��C�|bW9��D�٘/r%U<Gg5��F$n8�O4U!\a���ha����V��ɷ��� z���c�:��#�%��.ؓ�e_;�c`
��t1�����\Z�-����/����<$*7�_���g�H�t�躨Ȫ�>�^_��F��ݢw�����O��*��R#��G�G͂��}ڄř߫+�Y��c<�Ml���2��ND�z�e+��N�؟u����%㇟���P8?}�����R?���@�׎�sv�1j����Q�<q��B�� jn����]�:��.�G7�@W�=��h�-����\�\���<$��mB>��s��h�|���+�f���uD���+�Eb^��bj��{!�b�\$ǲ :f��s&���͢-%���~�H�d���P�U�t�SO{�G�������tm�5rO7��j�4>/i���]�0���Oښѿ��R�Y�m\�E�ϭ2�;�Rw��ں�(�� �_�Q�v��M���t��_�4{:��ܼ���O0����>��o��&�<����t���/����k,FrT3DI�N� k���6�o{��Mj�?��؍m�$�x$������D��+<�d՘v�)� ���>��!�7#����c�ߵ�z��E�Ѐ�jN�-=D\�u���'/%���yVҶB)C�ӺUW?Frߐ�ICu�cC����>�&bS�W'����������Q�,]@�Bp�W2�T�韆#���|*�zV�"fZ-�*�/��u!@��֓��B�
�N���-��e�BH���#�h�-'T_�,>|�"��U�W��\���
��O����|/r��f������~��)�J��o�@k��&k����Dj�����PR
�켁nq����J�DVs��~��gL�����1���Y�P�0ֻ��W`������{**?	�ɼ߂?�Y�.�[�%�� ��Z0r�-�~����#�w��瞯�D�
���j�⍭������J�3�x��u���|�_�uF�P�M�] w6�Hh�2	�Y5"��ߕ�����g(SG�]�l�$H�_F��ϭD�Ių��W$с d��2ub;Qݫ����� ����L�b磖�����g�vG�D�BS�G�s5�dɈ �Ka���F,Y�ʙ��&rH��v��s���!��k��$M����3�mE���C�gmR�EA������ �}�>�t��q�_4:� !w��ΗbPf&��AW����غ^T���9�hTP�y+X?pP�Xc��f�^ʧ�xk��7uw{��ݙF=��4.0�����>���CY�s�g~9QX�����p���x�/�#��A�z�N�:ې�f���KQL^�y��񁱛Gc`��t�u�JNim|F��ܕ�a��� 舊������DLp��o������e�X;D�$���kG�
pd~0'���ѷ[��$=�!cs��eG��ck�nn�N1�E!�$��a�}
t�>!�.�JV���YNs�R�ߐ����"��-K������ 
����Ѭ�[��;W�M���XM�� ��D�v뜰� A����mSzk�I@>Y�}]#�'�yiY�j!��4��<�����X��i���GFM���1!���X �XU��2A����p� ��p�[��^cU}��\3?�7�ʥ��˦��~���c�Ղc�|H0��D:�~��� ;S+�9g2��z�wB�6v�q[U7�KV�e[�<�hg~h�b�\H��Q9� x	�� {�>�_�P�(����Sɱ=��w=,,�_-� �"ߣ���MS�~�ů	�6	hz�X�Գ�3��N��2�[��Vۧ���O��b���N\:�j_��b$8�B��5W��I�z{��HR,Y���f�o�ER\�¬���7��fp�|��,Ž�|�r�[�V9��ɶ�o��٢̫.z�(��b��|b9]ݚG���9(��(����KG[EՓ�$$�sx_��ǟ�,�������I� ��ơ�{>���	����r�p�@z�>��Y�&��Ǎ���6�N����j8��q�������#�-�~X��3�I��oAr�I�RA�!��Q�e�jV���aP���.7��to�gH F�`�GBin�+�+Wh8�������{�Ѫ]�V��fTK��\A.|h�0:�b���"�w�j�;S�Z��+�j��xg
��������M.H	�sGdpF����������U�p�es㧰���d�����!�
\5�W�Q�u[xb7��X��%W�o�ga�H!)�.�F�G���T���1�;cT��z��U;*�n��ٙ�K,�'ƕ-�%/ؐ�����/=�E���	�ɘZ�7�3"�@O�3�[���^Z��C�p�Vd�[��mLf*�iU�U{�p��׌"#�f�f�y����������Ĳ-fu>�$h��|��@�pZ'�Zk'0��"e�2B�Wm[6h��ΐ�P�,Nd�c�0&ߵ.���F��8�U�~�%+�0�d$���쁂���C��5��Q�y0�8\Ń_�N��ݸ��������k�)�]���(ݺ_��s�^j�HA�(o���>�����Sh�y`R6l�7�6���iw����C,
F|2�/�;�{�(>-h�v�P�5����α��,㵒N^����^�,��s�sͦ�Я��5�pu�WsQ>R�CYk%M6�͓��L���}˽Զ�a�,�m:a��Aup��tV�v)���U����4�^J�sz�ي^Gͳ%ެ��0�Gam�I��6/���i9rj�9����R���-I�J,��3����ܮ�Xv����X%�+�퉔���3�' ��:^��<� w�?ӂ3�Q��`�[�J ��w,m>��^V#K����3�9K�����ǻ�ښ��Ա�!����u�?t���[2+�<w�Se7���H�2%ªhf��D�p3�"�w���.�5��O�����d�S/_gم�T6^���\�'�]n��_.lzm���}Ƅ�kc���=�Jwy:h/~�p�rw�w6w����׭\��W$�d�ba4aъ��xl��㸝��=��O��?p2ʢ�}���@;����(*��4��"����F�YLE�X��I�|�haF�#��aJ���lF�b�ZWYbp�v����%���M�A�'�=l�."j�o ��h�8���H�@���Yݱ������s�_'��Vq��A�͞�"9�O�?�)l�
VS���q(,{���Ѳ פv�4�зܲ�Zm��S2�0�W?Z�������J.�QCZ��Io�Hż����>�̝i)�M�'��rD�4�� �\�r�*�h)}	�%���\u���H;���0�6T��w�Z/f�� g�Y��J627�&[c�q=ʭ��ɋu��Y�:\��ݶ)0�����,$mr~{����uh�(KϞ/����3�ɳA���Ꮇ�A0~��`��o��4����'ZN��1�J�u[�h��J��:[�ĸ숽�7��)yVa��r~�z�Y���z]�O��ڢ�:N�G�Rk�5�7����x�ж�j!X g�K�����c_�д��x�V�u����Ʀ�Z-`T���kaB���x��E����|�}�I���Y�޲Rw�f?v��W�Ɍo���%��B���U5�ׅ��ul7ZO�Y����¤2}vh`qL��9��"���U�'>�w_1<�ԩv̢������0<�AbD��x�����TLzR�N�dY+�����_ζ5uu��dw�#3=�s�^.ԓ���򍻖q�l#L��{��*S�Q�=���A*<�)��
��p���orw�Nx�q������Sį�?X�W���|O����2�G��~�T��]��/����
��-Y���h��jD�}=;;���lW�^�q+P�R�����@�6Ժ�3���}X>{��8b�z�B����'OS�t�9�]���i�_�t��,����WwN��й�Q,����6���|®�W��2E�`w�P��>D�=�%�6jH����R����L��U#��H%���Y>ŧ���	/Ҟ���_�?���W")@ÁyQ7�[��"���Q��������u��/�a$�DD=�O�E^�s��fŤ��3m�A'��yo�3����>�sT��g��rQ��1,]���b%'��H;"�i ��"�'(��j�\9�������^�J�^^~�1���"��`+�c�2&;��טǭ��r3������<V��pV�"(��}c���(a��H��Pg-e �9Ӄ�
")��."*T^WuJ��IПx�n��S�J	39B#�i4@bN���FT����X��K�^a!�I���ᩨ��Vy��7���t:��fb�'���߶��}#���5a��j�"�3<:>��Y�ʋ]�
r텴N�8*<���=��_�F����ݞ��ɓy��g��%�:��5�Q���ߝЙ�����N���^Scp��I���~V�*�W*`ӋrL����237fuh���c%Z�&���N�!��R��!8���M�>$ean�o��+����Z&�kN�}���0�ٗ��L�������}�M������h���]��u���X
����jE���m�2Bܛ���(|���o�����R���E��'�H�3��� �on�� 7�M��^�Y��^�Nv��=j�7V��	6Ɉu�W���]Z�(*s}��I7����d`*g��Gm�����Cj��3F_�Gw���t�V5{v*�s2�&��.k���o�z���`�����RB��w�&�������|b�(R�iJ�z�&��7'�Ul0"-<p2�M{�._�&g��\ʧS��d[S���@zCS8���kaĔ�xT{����@�v�i3�H_]d��v���ˢ�pe������Y`��(���'&0���kp� P��
ʇ�	����`x��rH�4H����ɶǯ<�f\�)yb�Ru��2h7��S2�\�	���s�� ��}��cJ�_ ު��,XB��N��͈6s ��t$��|�B���M�Z��lFR��Y�f8���`{n�n1���`��EK\[BR���)*ay�HHC�~�� �I�Ƶ6��5�!��2<Qϱ�P^\��[v�r�����\=��K�k�M����W?�Ă����%��Q���GX猐6�Ҙs?�p���E�쬡>'@0�T�r���D~����aέna�͑y�����k�s�&��D!|���FȈX�� pt��` /Rn�=|�]u�в�;+�TLt���=rㅟZ�&�豧nDg�e��ϖ�N��ik)'���/EvoQ�Oѵm ��V�qt v�[��8�i�ۄ�*��4�[@�������ڹg���>��CAu4�e����ޙ�d�؂����sիx�!w0C�!��e�v���[)������a(U��Ҝ��),"f� V������0Ⱥ4��.jy���R4�P�;g����ͯ�%,�r���b �bC�}��Y��F~V����Q��N���w�����K���"o�v�����6�~{�9���	�f�XD��:|��<�P)ڧ�z@H��\�Y�T����G9I�S��==Q�>��D~��㛫�Z���wk.�g�ћ§����d6���!�/�l��=v�ȯ��#$|dK���T��CG�5s��`@�d�m��$�M�u:�O�Vá�^F:�XC
a�׺L�m��u�T�%t���q�ٔ��~����]��֙��i�p��"��ڐ(�-y`x'%m?�\9��8��/,&�e��ɔ>W��y�������A�(L�'J[����>���/`�zt,���%e���W��9ŗ���=t5'�s믏�E�q%zJ��aZd�>��G� M2�	�6�{2���h��֩Z�k��o��׆��7cI �� t5���U�jj�c�ȥ�0�]8r�Z�|^*�r��߲�y�$Wz��#�Y���ċ������"��'B�P}�)��l��:񮯩)�r�����ި��@�MRa:ψL?������^RIY<E-��j�K������sHB�5+¦S���B��Lڀ�ŉ��� ���<b�4�6�jWd?��*�'�tI{	�~�2����+W�;VG��B��xS��N�KT��\8}�|����@�ɾG�<��ہ�!�@���8����i��u������7y�*�NBS,d��%�����H���r�=��^�h:ͽ*����q+�`V�8Kl��e�E�8#���T�uvC��!��G�#�K�+�h���M%f�P�D٪�dNN=�K�I�U�~����^W.�%H:0� F�>�1Bf8�L -MP[�D+aA�B���sV��a�C�V��d�1�D��7ݱ*N�o��8V^	��a�/�D�e��Ɓ�H(�$aaC��ϒ��s�nK�w�(Ɋ����M*�8o�y<l~H?(��	�oT��L�u�7^L������+�]/�VW6�o�ґ��h��h�����4L\����/o�s����ga�Ӑ~�o�Hc���b���p�#��'c����
${�݋�l�%�_���+Y��a��_4'�%���q4����ߵ �U�=� �WfQ�+��*��523 ��x��pBv��h�����ݜ�&��|�>��x'
���%W�[=ݏç9���.b|͊�e���_D��.Ӽ�ȅxn�4͝�����K��}��7���o#��P��@U�X	=8��rv��&�sW�y�,R}���w�Q�u�'�jh�3z�{�P{��'QD��WC5VNzp��p��L��]8�(�+Qq9��ߠ���/��N(ޅ�o����ibdW�)��F.8"d(�Ǽ��@jUt8����|F�f�打��Yu���h��C�ܗ�.�l�"$�%~4Ō٣�J�\�P�,5�i�Zb؋P*�(@XF�:��6^Mk�X��
L��]tθ�&��zm2��D��/"H����N�R��B��n��dz��r� N�R��Ǆ9�Q'|�>�y���>(1�";T`��s��B���E@�El�@ p���G��ʷc��5E�9vo�����{���a~�1y��oIsF�f%���\o��|�0���-��:�n�|��,J�N�8�q�
��6�hڇ@�'p>�~��:Іs"�hb?����ĎE��ݍ��u�h� �_���'�'�F�b�Q��p�o�X:��.��:j��K�����٢&}�)y��̎,lTLCþT9H�[s�󇋆e��,��Pz�h���-B�n2�u}e!����4�z�7b��օ����+Ħ�E�FG^�K�O����Ы�C��.�[�������%3�uB��[p�UqؘB{�A�l����#�(ſ-�^��8�Ej3T` �y0*�>���@��F��-��Fܺ��H{�Z!e'���*��v+8"[�����'�1�ֱ~�L�eP<��tOX*��;��T�w�̑�1�WZm��C���y��iy1Zi�N??"�>���Rr7�ּ�<�Ná���� 2������)�U�@g����������}�<��s���8+YWU����F��-�ı�N����9�!e������@��QC���br���K�ϻJJL���y���x��ќ;ɩ�6�SSfKM2���(��~D���ǒ�A��rH�R!��R���Z��
N,��.�j\������o�㹛�Q��;��$�&�z�]<�2feb�4��N7Y��h[����T��=$��5��
��k/A0�Y�E�� �Na@_Wim���&�S�E��4�3J}��5T�u�"0�]%��n�$�����q0UT]��P��4�0��E\Pp*���(A*�H�\>�o���ֿ��#���˝������_'����D[ۃi�����`Ԑ`(GM���f#����*J��YW�����'��)7d���z�f�П�9�.f��~�:�1��Ǘ�U�rJG���CcJ���,f�L(ȸE����`i��9�'���bT�	&�5��{"P�:�����&�e
[?��!<���6��R��:6Z^���_��ؘU7z��W2���dIF֩E�lFѦ���C�&/۲��
9q���t��DP���wP���T�޷����a2J}��:�/z�j,¯��%�:��V�,\iQ�vKb&�N܄M�g��p��#2Z�Ķ?��O���>>����rȈ�!���|�`�%Wy�����Td��+���	t�8���`��j�ş�����kk��� 	kz��ҙq){����į�5�g�{)r��
˅j�3�	�S/�g�nv5�/�rGm�T���w|c�dF_�t�m13�A�g�(CP 7�"]�9�f�G��(�BP�Ŝ��p�����[0UY���l��r�ꌁ|�zXDrf�؀u1z����n5��6�����\^2���5Tx��Y��P��d���N7���V�F.��{Q+kaSfv�� �7�5��U5๝�	�Yd'2��|�;���+�n�,q�+5�6Mt�c�Թ� �A�}t�!� 6�������H��׳2q1�v���T�ѭ��X���;j��z� :-�v��xy��(�a��~��{3���W7�r�a�@�����*���|;��M��m��#�&V���� �䑠��!�	�f4��b,"Ū�V]��㔟�G�W
�KJ� ���|
�B��(ЯZ�B��&��>%��-�|���R�=º�o���Z�����ܧg�G2�L�v�q�*��w����_�!��9�H��<={�l� ��k⪔�)��.RB��P�fw��ܶ��
3V̪� �{���PFS�v��2���xEGH��O�9}UMQ1�g�A����i*��ɏ�����<��U�n_��$�J�^�+J�|�,�o4^Gd@l4�أ���.������2������CF'���rH�U�`�`��#��]�|�r^���A�tۿ��-ަ9	]��x��ft7�'b�B��/χ������		��2:}�kQz�iJA=(�����57���dP���4�ނ���>����
�N�v))�~�U����i�LFE��i�~Y���iv&Y9���L�#G�8���,�e%�J��V!���v~������t��0�������V�G@�p��D��T���@?�ʯ.*�E��g���\e_�h��H�~�(x�X_�X��B`H��U��������~������E�?Be.ǻ"��Չ�`T�H�
s����(\�CV�ڸ��˃�q��;�G��N�*��G��D���U�R��qm��Ƞc<��Q�f��_i#x�e����3���3r"1|�:���E�8l)��.�HD=�IYx��,;�#�o��;�N i�mh*�}�4>�	�x����9^��/�|�R,�K����ȼ�̈ǋ+��e;�����]�~Y�;��� X�=Ɣ��� x�&����	/�q	�U�����f`[),�hT<�ge�L����1$B���)&��d����6R�͹Ӯ�ܕ{؈"L�u�~���X��YyU�
��z��3�c�Y����:�Ք3e���V�0ڶ?����~3���l���̌�S� j1d�/U��1�����������wv�G'���/�e���1��":y �@�ɫ���ϯ&�6�פ���Wއ��͵Z����y{p��W.X����Tݐ �XF��@��ƍ�|
��YO^oE��O���O�YҺ��!� oe=�PX����iUԬz�]a��,� ��ල�]�݀MTڜx>�O�ص?	��C�=�jb���>�>�"m�A~��F�A���1����î L"�����!��n��,����=�ƅj2�A��`7@��O�j�{wk�d���<=����Q �䱌��\|u���4�~ciw��"��}��,M��@��g�,ynl��k�+�ꨛ:ɉ��������NVS,𘌾bt���������aAW�E��Z!|�=F�	^�Ѡ�h�1�|5�_b�&��Q����m��7����Y�`>P����uIw�dD�Y��qA@�^�s���(9�P�cSK���m�&�$���AԊ�J9��X�e#N�i���5�M�!#� зy�C�"µ���_����C��h���o����0M`_zt����5l�J��^��;$�� �C��8�Cý̂|0���6/8t'/��&�|:�n���6-��^��9@,h��e��rL���kG0Y���Q���"G����>��Q���|�:�����-iY4����U�J�jY8�,wm���S'Uk������E����]�&�	�V�h��d:��A6�kP�ӘdT��z��I|���|����ȗ��ל)ѐي\[�[�N�7��!^�Љb[Y�i�QgO:TNZ?�Cc��P�b25��r���J\*ndtMK�h�#ٍ?P��v[�֥���
�'S.[æ�怾ś�[��� M�R�pLcƜ�O�b��xzG�8�qc�v��p��ȏ&,[�N15��7�g�a�O�����b�,b�������-�Q:�J�S�<�\��n7L���!5�yz�����f��6�Gd��l|�"�~C�hV�T�ͣ��r��n\}�n�������
\n00s*�J�a��{D����/a���r�%-�^Ƃ�����9G�6��K�=(�z�*���
o�%'�B�B�4kf�G�Dۿֽ�}b�a��]F%as6
���x/���a�����Ѐ���j���W��X��u$�KD������sK�^q��1���[�e'�"�Q����U�|��*HA# @��\�k�4��l��O�*u&�+-�51h���`A�N#L���.u��u��Y�#3n�*n���&xI���Ywaщ�b
c)rx��%�"����z
��$�q��tbR�rF|���̛;�Q8Q�xeZ��������x�pX^�,_�~.�u���9���	KG�af�D��n�]=�z�֊J����}�/�N$���������g�V�P`���N�Dfi���rof^EW+ڀ��Le�Wag��'�	Ej��:ָ�N��)�D��^-����shcϏ>
{�էh9�zg�`��pz�n�mG�q>$Aԏ�L�[��7U;��ARo�����H�Vf�YF�ϙJ���O�Fz���'��3S�I��SG�Ɩ�f��p�*�LNR� ��d��pN�c���P��������:V�k�.-킲��hG�g��2Mx�y�6��q0Ϯ�����l�`H!�GX/�t�,N�E�<�:��9�ԝ��mZ[�ƈ�:I�Ⱥ�5R�R`Ɵ2ÕB~y��C<ݰ���2�!^!A^r��R W�$��)����oM�`K�h�R���|Fe%�%�g=�;B�;����r�h�{�cN�N*V�o�%�k��fo(6�A�f���9�٦�3,��\��6�}��}��^���r@��QUJ���W��ؕ\���_Om����Hx[�;%�a���cA�bɘ���C�@������w.�b;i�bg���ּ�+_j2-#+��J�9�^Lʍ�:�*V�.������Z a�,��7M�u|TM���i8*]�J�'����-ౝ���T�j奒PJ��XZK�o)tZ>��ݍ�� x�d��k�����A�V�C��:�gg�YU��m0C�_��wS~������C�P���7��;U��ܟ�v�&oc�g�@�t���k�C^GC�VZF�����~���aN�`�P��Y{�O.��R@�66����{�������`�z[�r'e�Y�GX��s�C�Β���p{3t�D�
��Il��wIN�ךO���+��s���/��.:��Y�WdR����<�C���/b �Y������y����j�QF�3hYQ�Qc��'���p	� ǂ����sDF��;����.��'%Of�@�kp	��/�.��'Y���@�EP�� e�;��Kd|[��g��;����t�ll���#��^���uU�؉ck:�<�6�&��F�P�pM��_M��ޝ���~]��v�7!�����:J)n�b�u�v�<�W��D���{��X騘M��]�.W��L.ֻ�W�m�-_�XaB����(h�u����Qv�⑈�l�"����H�j�>�E�9tт~I���ny�'�x��yI�N��4*쬁��?.�d/�c��gp5.�B�_2	�����YE7�������r�\x�;K"��Wڧ�F�q< �� ����C>Z}�=D�s�x0�t�����w�a��1���)�������޿+D-�c��R/�;J ���?A��=_N`�����H	�υҺ����WW��~�3#��Y��^η4WA�-�@3���B���Q��f������^�CA�(}k{F5(ߧ�aK H�6�P9Q�li��������"I��a-_�,}݅��YA���k�crwɽߞ^u��1O@0�p6��dom����WR��V�m�̵�\���y7v���y��@ҥ�lg�W&<]�|h
���wRİ�&:�����5Y�x*�K��yE�8�x���]�i��ֱ���]az@z��c�Ir?j�8��/��ʓZ[I�������#�E�����sQa\^h�Y*C�3�����g�-�;�vX����)�F���K���V|t�7��3�C��~/L�F�,��C��� ���ܙ�r<��<*u�9|�����,�z��=�"T�Y���	�a|_�J�Q�D�Ğ^�*�rP�9i��d`����a��*�/����W�oi"~�BRo�����:��X�%�������Yi��Q[���u��Б�F�n��詹�=��o��v��$=1o�=�I��3�e������lo�8��p�؛p��V����$*�6G�%{l� <��~V�>4:`}���*��?g�ov��� ����Ȥ� �� ���Κ�h�)͋��ٴ��&V�'��fl�>Rfx��3R��<mhCr;M���!ớ�'6ĥ0Є�FN�B�'�]���+(����̏冤%�	�!�q�ƀ�ȩg��@w �Zj7z���'�Y�bjΝ��!�,$�����	85,��5'�$˔z*3X�A�Fi�����
��V���H�71]�Yn�kK�m���w��Ps�3ʣٌo�G�<�de��S�ɰ��?�ҏ�Nn�_�R�t�x����JxVk������T`���N�5���̋�VYE����0�c}�/��־�鐤?�jTW�+�wG��.Qp{��X�)͒K�N�/=�����֫/��_�kZy�~�?3��'hE�W��GK�.��<YD�4�b ��|:�&����F����2�����ʣ�Eͳ��QD{�.�G����MO|��i�x	�mίm��~�:-��%ϙ���$j]�XK���|�y��g�{�y��}u�ݓ��?R@�2��`�?wG��O+��>�I��}r�uvU�g � ۗ�׽�(y`-�]A�a/;��g8��6���O��}���G@ӆ�:��С�t��]�X�4#٧���Ni��Q楿U�r[��s��}��Λ�:���M?�����\��"imZ�.5I���?�ѷg���dR{��NX�����S��']�7�2o�vV&�*P�r���e������Q.V�1���Dw��64����0o��Nq�s����>�?��_�ZT��c��Ʉ~^�њ�G{�͹I�*=v�P�4<��wk��²�t�bG�2 fR)�'����w���&Va���״
�F���7^ �Ą��;�d~d��Î���-�����	Kg��N�=�;V�r�J���8������֊8�9��re߅r�)?�4���m���e�*��2([��Ȝ*�۷R����=YH��ƚ����5T�Y6:�Y�_���WOR;_ꂬ�L(�&&uE��,��-�x�v�3���l��y���k(f�f�i������"H�9��_J�����J_D�6Җ�O���W�Xg͍.9V�o�g(�e*2���QT~��iXu)^�����S��q}sl�$Gns��X �4�#�F�T��jf8�`{f��`d��~���T�`��)�>�6�M�G+Psバ�i�m
�A��>}ۊ�%�~�7v�Ը��Y�"KG�:�	�yK�!]G���Q��с�5��x�se��P�?�s<a��Mj3$v�+�L|,�З�E�/��/��Y�i�6uz�)�D!j<+���v������7�q�p�[����/hjR��.��#g�����9��?�Z���hv5Gb��	���8�9����!f�L����K��	������?�؇�Gˑx-�}{zR��t	5:���_9r���m���a�cP�syx�m-�D!rl��v��ۏe��ЇQ�0C�����cp�P��
�֣��o�����ֵ1���Y5�YO���![��,a�.���8[l�H�Ӣ��n��R�:����r'@&#�Zj9����xخ����ϼ�0#��ɗ�1��Qh᠈�Ƃ�/㍸��S$݁B,��0�ʝ��bȱo�Ҳ�ܖ����V����56~bj�X.���������L�![t~� @��`�Q�rv����U8�ɚr��J�vZ)�o~��[��@�y�N�`z�q�Q���E}������ `aO�B����>E5�HT������l5.T3��>uъ��f��^�⭵�{�����x�I#���e�$0W�r�
3�[�h^8a�h�;�^���U�Aܓ�q�
n^
��b��)��т�r���r��nIEX���"�8�5�z��/����=��3����rhH:�h;���׫o.٭,c��8�:dC,���c\̬�"w59�|�T�jw�n	�Et��?	(��:�֔����^�V�����{��`x�$׬&6�l�h�`�� ��+�퀚����;�΄�AY���y�C��̴c������V��wp�JgX���r�//&,M�~T �/�HMqQ�$�f3�u]�Y����Ej�H���Ȱ��"¨�l:��*�Y;䅃�z��>��1J�W<:����@���r��΄�`�����c�;v�-8�b!�r��w(uI���ϭ]��坼'*(B��#x���ޅ�ճ�Sny#�`fn�R��,ਤh���򭌸�����mV��8+�[����9�ܐ����Vg�K:�_V�9��� �X_@s�v�׶4�_�E�ו�C�]���O_det?,9��G�ǣ��	������Y�@�2T�KbMF],Dp;�a�~�s��@�U ��g� r���_��Q
+���	l�b��Wܹ�'��P�uI��H;QQ��C���i舊�'���1(e�q�T��$%j���t�fS]4X<�م>�.c��+���^�N��7�_�wĀ�ߛq-�.��x�~�`@���F��$�1�*a��jfc��p6�ZFk��8q-��9A纈����dwT�>���Y��f�{�MIo8])ލ�e�2�*���Y����׮��䮝��"�;�h�8v7O��mе����c���y�,p�%ސ���H�Gէ���%�P�Wq|���ק��`�x'{���{ᬓ�ˍ���
$���P��8���acIN�w��NZ���/b÷�;�ǏC��i;3���^U�қ!J�3jʙ�$XH���s��9�}���
w������C0i��=k3|���H���z&#1tI
Q�S}�6O`�49A	�}]������>�ڮ �����Cs�Yh KƵ	yN.b+��e ��z�O�X�|���$5����t����z�{f᫠t��H�x�������/�J~���M�y�z�d��R9��w~��2D���:�
���>9����ٜ�ER�z%�5�T}ǟ�D�_�{�o�I*�EfE���^��<��}i�b���'R��"6��O/R!�� ����� �A�m�n������5�e�^B�� �������4<'��-�c��fm\V-(��w����7	�d�c�p�#y1&.u��,%�4)j�횭~�@_g�K��rm�a�T{��f<Hk�ʯ@Gs��:�=���7����aſ�:�s<m�c��-��� -n�8�g�=�_TO��1�� K_c��G�Ԙ"�iqB���E�O��2���C���"��{<Z�<y�p/����M ���N&���ۺ'�jnL�m`�PLڤ0�#AC;��]*�H�caL>-(��Eи�B��t$rSP\���a;���#�2rF'w*����$�H�I�ʧ)%b0C��?
��i}O?隷|Ԫfm��?��Ѷ(u���7�����Ce�B��ϠZ�ع���Cx;U36��!{Q���EJ���g7�����H��t��:'a���MM�HZ�5X�p��1Ŵ�#`�S�7��;ݥ�np;�@�b���C$���X�������m�n|ɩ�,�7��J;�*>��Vd8,�YUd�`��̒����[˟���^�aK6>�NfT<��J�n�4ϵuN�Ѕa�1©�:��WhVk�#x�H��ؗ�lO�����_��!�#O^.Y�ٍ�`�"W�"V��Z�~d�EC�4�-U"�����,[�%+��sfڋ���˃5�QC�4܄`}��\�x4ǌ[�@�#b�zZ]�샎��k%�l����^S�+. ����m�ή�Z�%��0��|E̖��^#���w�wh���܏dH�9i��{60�K�R��	�B�!�	r� �IsV����:*��jL��ѵ�d�0O�9#tm�b��U�"���U�&�Ԁ~�wk�����X?C����hwζ�����Ю��([��gh���ᳯ:��@���EH�7����p�̮���>�}��g����g�{0E�}`��r�Ɋ����+�{-��M�>ǋ	�UQ,a��a���d��L��0�r��q�-rR�B���pW��)�%T���v
(���]@���<�t�6s�en����$�l��W������i�hj���[Q�ד�� �-	�m�?oұ��#�t]��o�����J�7��B'1\�߄�l�ac�I�6��-�+��t���07�k����s�U-b��ė���Q[K|��|���l���q�k˓6c�}��y"���7�/A"'>(�Yx��@�As���P���;S��� ��fLY�	Gġ�>a�c��	���3Ñ8FQ1��@{�C���2�@��*e܏�o�m�XQ�ʟ��mk�'F��
�%	�ս�<uI@/$�Sѩ�S����<����q���,�ܧ���=�7Sn�7o@%À:��o��f���z���t�B̦y]a#9��)�;EA�a����}�oL�U��8Z|��IA���XNe㑥7�� v�I]s7�O躻-���E�T^��X�3��T�#���e�)n_�n��)[­Oym�+,1Z�C9bi�	mKlA�ލ�0a΁� �D$~7��ʒ<��*���IO��¹	3}�V�>r�;��=X��l�k��UO8��ߔm�������QEL�bEv�� N�n^g\(Ǣ��Y󮻳����J�\��g�v�.˩�]�&%dhn`}ZM��P~�lHu;�"s� �q�%���U�ʾ��DLC`���C����վ�|�-�U��q�B�Q�hq3������	�u�ZM�8�:¬�φ;��݊
|y�%c�pOɠ�)[u�6�66���z~�>J-b�*c40�Oِ҈K��#ך�w�l�<�R�v&;�e�����	B��6�FZ{��]Kh`Pw��N�*��l��8U�Tpw,�k>'j��N������n�v����W/���Mq��<|�&yZ����_ٺP�+�d�fhrȲ���4^rb�([L��:X�
�·9�5���l�~��ڬk�E��)	fG��
̒���6��TK�t�>L+��[�7i�!�
��$%ϫ�������R
&PT9p���/���xi2�����dȬۢ�7�9?�R"1ƒ�=H���WK�fNcT�q�5
��Ą�
�樝���<�@��/��1�p\�#@�#e���+���j�*��!���$�C��&W�4tr%I��O���*L���>^N8�+��P��ƿxPb�(�3o�p+�u���ᚸ���Ґ����*!N��_h4?7�,�Kz��B���z��v��g}+�Ȱ���"T�L�$�x*�}b-���;5=eo�ɤ��G (�r�~h]�l��="�vP���9��Pw9�W�J��mi-��x�gc�'3Z}}����\�1h �R`��?:�o����5��es��h:m��4L��}�xgYH�/#1�����M��*Q-���X+;V�=�O#�
�E״��#��&�y��vH���%(d;/ ��Le���@G� ���ﳾ����d�|�2Bs���
�Uaj����%Id:4:ρ���EK���7!eV�$U��z�^��]����ۀ6�\�<>�{dc}xf�X�ɣB� ��0�Q�����s��c嚂h�;�Q��� °���y,{���3����Nl��5ZB�,V��cȶ�'�>�#vo�o�1��<
�]��V�8"�k�;h`��E�B�������΍��t_�n!��.��w1�/�3��l/�SmM�zR�K g�ruϚ�:�{���*3�%b�CT�_@���X6̳=��p�k.��͐��}'V�Φҏ�i��4Ok�n\�n�y����ѯ]����!Ds$�����v ��>G�]�8�W�����Ŗ��!f�G4�S����=�7�N6� �`��P���O+t{��Tstȹ ���5X���ߟ<�lX|�ƽg�"��a�O��+����{���*���-�R�s*������=�h���!����`s�%t'FI���>��<͍��)�����[���XUQ�sG�-�(z�����tG]4v'B�^��Xg����Ț4�	#�.����R�	�~���,7�hV�lQ��x� �T�S/�>�WWJt���
(�,�G��2���7kQ�a�F�;��!Kb�xU�U)��3�p�:��G�]�eF�������,��=����r��L��mټ �������(���ܷ��Y�I��7"�� �P�G�m�6"aU00��'���+ؔM���Ls�z�bǿ��>�e� t0��_�d���0a������!'n=�0|ͣIC7Ah��YM�b����x��k�����,��i�UvڌM�����U}��p���&�+b�g����Ĝ���dg���ȡ|��pW�:�7����=k��w�"�yf
�JI#�Dz�#r��ʬ�o8y�\��۔�gics��Q���d1ҙ�KUw�v+���t#fR��<�X���;+����R����z�v�8�7�A�9�"���zO�"=�&^��Iin�J,M�+SD��61+�҃	|l���J8/P�"����l.oG^J���pSX4wV��~��ސ�������(7�Ts(p�e�+d���6�.@��ێ
�qք	�����	��zן��h�?B�D����̕i"<&|j�E��H0"�����zr�ܷ��2���N�!:C���D/ ބ�)��Li�SԀ(>T�RL?�T?38�1�6�	�I<���|�Z���7���<�J�~�~J��J�|W��Z��{&����-���&�MI�JW_�W֎Kh���S�y_D�3����?k���EP�N���e]��kb���l#�C�U������Z����z�x"��I���<�Y2ߢ���G�=���^�U���Cs����,/�;�BPB�g��{��p'��)���F�g����;IKL���<�>;I负d�]�Jg��5�CN����VF�q\{����b��h��{!��[�v�e����^L��՝2RE1��3$;z����v�x�xYK�M,���C�3τ߄����	����r��u�������6�;��J���eӯIGUy������-�Q���ԁ�d�am�!��C��/�`�C�J�ǟ~ �i&�Sw�;PTA�J��w�T�4����u��*�!���L�|�Ƨ2�V纯k^aM
-��x��J��nw�β#�鲳�##��W xpS׷~D�Ej���-����EA(���b~ �m#�/�0g�yg>�� �E��h�;���᝴|t:K�+��?/�B��b��1�}B��*���cJJ�B�;]I�/bD�_�ƓC27|�8�P�������b�,;.̘��>s�0&���5�ff�y��ں*�w�Z��%Y�/��Y(�>�n���W��!�z5����|)���gRT�~� �����o�do�z���bNQݗNC8Uq�'I��E�bW�v��	�e1�dcݥ�{)&l�	�v��!0:�0 ���̉}/�m��Sm��!P!`-Gb��>�5�|
f�d�����Tb�^��
 �lI���ew~-4�\�Y����8.���G��ϯPG��r��DH8B�������2�V�)`�/r\e��?0�E�\b[��*%w��AWNF3�%�␈El*��>��n��킮���mo:� ���ښ(�������[z%,*,K%v�>%�����w*�8��᤻����V�pq���Z��Л;���82r_E6��Zb&�O+f[
܌$��솧f�����N��>�R���!�b���p�9?��z١B��T��E�)l�&� ��� ���k����Q9���ȭ�n�H	\j>�{%DT�P��eZ�4����A}��}ilR�O�j-C��z9Р c�����^��/�J��J�?RV��Ja#��2�����$+��Ck0:|sdǤ�7���G8r�1��r3:�V��l�~H���s�Q��8)9��Uar�P�A|5��s�J#��&z@����=̔��
�hȄ��D0^��彪MU�?!7̱��7����N
��x}�5�ٓ;�D�]S�ښ�o���#����, �JC�����[�yW˽~GPz3��}���:��fS��Ahu�������j���ւY���_��ifu��ltR����o�b&E����a+��T���~hC��	���6���>���?�S�>!�l���Ɗ.y2H�����Ycx���=le5~���n���#���>��\i}�ڒ͓��P!��fb����˕-#��.�4����*�n�Z�X(ܐ�W��a�n���z�O_G6h䲭�h����A�kAEb�͸�pDq��H�����l��x�	{��|�a�?DH���R�/�c�"}\�N���-�O��CL�t� K�经
��d���C=�5�BLU�,`ȡZEg�E�v7�u_q��} ��R�<����	�ǃ�*�b�`:h��!�:X(�%��445��=/�[�=	~���+l���fk k�GS�tuV{��b'c���N�{S�F�+�N"��oRS�0|
Y�;�"x� ϗˁ�c�$�hYf}��ߵ�(ǧ�4D����RV
ɴ�/�!ǻy-t���ǣi�U�PT�xQ(�HFTԌR`enx!�E����Ѩ��Wt�t!2	�x\~�U|:E#Ӱ��)17���cݠ�[ 7g�-�Ȥ%��ʫ��jL��G���������?���"�:y�|�������V�W���"L�_�EFo � D��wL��Ί���ţ��L���9MTт �Е� �h㖩��e�=���S^�L_ڐi9�%��(n<��{���'{`Z��0����e
W��Gmy��Bz�Z6\�?���;����i�]Pu�Vr8�RI��^�J3������}�"�-���8��9;��J�C��m�+�7N�o�[���4��k�D���A�!�+����dJ�r�8���a�R�-����T�S�����m�2��`�h��O�� ��7D�eCM��⟬�.555MDǦ010��g2�$u�d�C���J���61{v�K�`�6�RM�9y�,�'���'R�p�;�b��93ixn5S�xd^��{�Y�Ƅ���"&�}�GK놉t��TtEQ����vІǪ�v���Ν�K����	)m�`��JH#������@#����V�J>�.am^�u**�r`�����TDk��lI �28
��W@,���#��a\yߐ��uAu�sC ��S �p�@9J�@0�m�`xA=a�b8�f+&�Z/
��*��\�̔�>)D��������q|�S�(P���/Y�I^������ӝ�8&�%��de�P��V�[v�{2��B�_ֵ��WR٭ $�'$��n�L���E�q��̴����Tt�B�OL����0��"���տ�Uv����^Tm��:�ޢ�粆�f"gR?�N�cQ*�c���i"�ꈦ^��������Ef�3��o�A�Ҫ�5�*��P7�C{ RxF5r�i��c�'�<�ŌJs�{L�S��!���KA�`�X3�kOe�u�)��uUѧi52	`=R��_�g{�K�lw����g��P>�YH@M�<Y�F+J���^�M��}vK�/΂vϯ� �ʞ ��,��-�hv�,��������a5��C�J%w�\O���}˔ll�����)��#�Ȇ�J���
)�%��%M�ל�������p:`�˟��O��P������U�Xw]P^��:3#k�&A�����(�MM��>-��aО��Q+�����+����I�V:�~��Fo��;j����ˇCb�^6z'p�f	��<:��U��!�����c���6��tʋ^?z�����ťJp��_J�C�D��cۤ��Y����ā/~oXLo>���)* b���#�����$���(�/e��[녾�)WQ3y�'��$�hL'�V6k�$eZ#zq���1]�A��/7����0@t���q��?*G�Y���re5�q��$�[/�ĺ���#2�/�j�	�o���Z��q�i/��x�+1�^�)!4�H�L\��6Vm^���0�i��dZ3��N!nyW����#����
m�i�J����,]!U���F ng!-��$D��m�U��Hf��v����FWJ_�M��z��iJ��Ͷ�����w|\O��Hd�̔���2����cZx4��i�.ߧ��\o�V�PW]�d�sV�qO+�AQ��4�<���MS�~X�������kP�o�(��M=�^f��k�·�S`���v��r�6O�h3:���a!�]���+o������(�����x��.��(�nn���ǩ�i!ȥ�'j��oL������{��'�w;����$��u��Y0Vn�l"0f(:W�q��M�Զ��Qn���t|�&��V@)��_'��k�2N�i�I�1��7%�VL��;������Y�N�f�cN�B�\����[,GY�.KZ2C!rF�-ٍ�_S˔M����b��$��(-���h^+:�-2�h5��-�t���̺�\yw��ھ����fQ��v�S��0�F3�����0��e��쩷r:�a�,�u�c3 o���	-"�97flcSJSJ+K��z��������z�����8K�ã�Q�a28/�~���IS�a%r��#n�U������]Le�>��Et�|7�(�g��s@< ��gO��d���+wZ����slC �'��K���mȘc�Zq��t�p�|~9�H+Km�lx������`}\b�������-�29@�2���ֲ��^���F#�Bj������,���K0@�h7Gޚ���X�FnL�J����<5�2Qi�3�<��#��PN�h �(n�g�-�jy��x�����Ѓ~�::����h��{�D����e��i��X�����y�'��kш��u�i��o�\6����W�:�[��'���u'5��2��Jg�u}�#�p����!�'e�4)�<Ĳ��*�(�B ��F9���1�k2���}x�*�~�K�N�{�]o�!j�Riw��ӭM�����U٣U=r��B���ވy&g�pȜ�9\���������*���p�/�`�!_Kq_[��e����?���M��VQ�fKs��*|�)��=��StN7��]���c2��˻o]n�M��qw\$�-G��(�1�o���w���a��6ݲ�vj��8�9=��J^(�ٱ�u`��	FC��)@��u� uW!:�<��u�WO���-��{[�.a�L#h�
m�%qƵ�7���⏧:�&j��K�"��C�r�/A�|��N)�& :�"��ɷ��6e͉&'�v@�@��ވ���]�jA}A��db���:=-�%��a���F����#��#o��.���o�?���o-IP�_�S7q�|m�iv�C�2U+1vN/��"Q�8=$��o�FF��h���ȍ@�``�\])SW�L�a�۽5��`{�:��K��WΤ�T��d��s&�Xm�7��#�9t���#��Q�F�G^���$ߺC}�[��▢����g�D���.Y��.j��������-��٠D���(S��$�fQz����f� ��v���+Qb~C(��#�G�2�B ����ܕp1F�H�vP/�6��y��B��fr�C��ք{�:œ]2�=�0��~��!t�g������/����~ ������x�aߟ��C�t���#�>�Qd`M��df��}�J�K�I�9����-r�k�
�MZ����h��5�4�>y��Gb�C]�]Ǵ�[���հ�yO�վks������b��R���'IT���߾s��@lI~�/��z��:�*�,s�>�D��nh��Y������i��X�t�6Cs���z�qClH)��S�w8i1Jc�U�ݎD��޽���%D ��sPv� ��J cH�Ei��B��"7%��YX�Y=� �U.=]��2<���եQ�k��N49ٗ��b���	�EkR��|~0�O�T�U�f�'�me���v����T(󲏝�p���ɝM`�iD��Q��FO��0b@�0��a�:l:���ǍER]L2x�����.}�e��6dd���h��l-�l�X4'yD8�Gz"�*��ϟ��A	����f֧gW[�;�����t��?�R�j�W˛��^�x.O��^�g�#_����S"�-�sͭa#K��]�a��v��"��}�byMq)b���}���!VUx�ݣ�Z�{;�� �)�"�<Y!�ƽ����i��BY34�����h~���2��֨�y�1���O �^�%��l�<��8�Ͷ�l���g�gV&�0�+���c>?J0�<�a^s@7�|ǗM���iV��?�������f�X�}����٣()������/}�o$��3�D��eI<0A��g�74"�ٙ��������K�z��9�ܡ���t��{�ܽ��64��ONN�-&��'���� Y*nކڕ�[Mt+!N�^~A�#������6���ƕ��F�_q:F5N����lN�X�Вr�~S������7ӧ��j��e�m@Ԣ/3?f��N ?�es�$Cy���I�bӻ���m��0�Id�2K����!�8&c���N|j�����{�C8�(ϻ
���ȴ!b�+��q����K���c�n�T����]��"��{�=}ƦG��_2T���[��}��7S�����:�ZFh�-@��,�N�{8b��P�:%�����H���0Ӑ���9��f
�ρ�S�3�o�ঁ*{ �=�x E��8}�Q]��W�#����m�5ވZ��+��S���$�s<��z��������Ĩ�0�Q#�Q5:�$C������L@n(�����s���v��K��j�����C�����0�ט�E��m@92�T�ooє��Ek�5b�w@�]��Z�;�"�jCo�6r%kY�	h��0�A�����x���n�s��+ߧ=A0���\�u�YXٛ8Q�\ဥ�V��6����3��mN+NQ��a/O��N ̡\z���}�x<�'7��9h̥[z�kR�#T���ݭ�HS��OO�$��jp��+ԕ�k�K�J2��#� )%WF�]¤ݍ�D���L�z��Uq!��]�;&�N�4T��l�M
I�������=Y4R��J��`��	���7�T2��� �Lbg⿍�>��]�g�׫ՆX�������!��Nek_�D6=]������F�]o"Q��k)�\ �:πO�peF�g�WoQ�>,7=��; �e��8Л��	� ��ܴ]e ��|C��u�f}������{P��y82���I|��yZ��9^)EO�iCT����
��"��+܀���r��BZ��<b��+B!;���m	d��ո�$=�s�����By�r+F��v���F&�u��f4�5A{��C��t��s6�����	[�;:�f�Y���O<��iTm��t�����n2��%�v��Z_���oU�p;I�#]!@Vvy�����2Aډu0=Kn�p�Є%��?���p��Do2���'�},���
+Ē��b�Vm�)�v#pA�t=�'�?��a~H�X1ޥ�����9pkf�W�(s��������M�	(w%��4޽[6Ip�z<sC�쫄&��G��&.<5���R��z�v/�Y��ΤYq�Z-�I�ܵAAX
MY>���o��7���K�g�`�2��?�!� Uzpܘ��E!|�g9S�@N�М��8��𰪂����'��i$@�Em�f�yi/K�y��EYIO���U�tn`
��x���Aԍ�ݷRgŰȘ���)��L��g[A���AO��eq ��("+�V������A����(GE����K����(�����]J�Z���4��Zx��?�]��ZX\�*�
�53�S�mO�3�V� �h�OVp�=!��(7����[E�����q���U����
 �"I��ߖ
 n�_�	�+dt-�,%����د*������R��U�?M-���CsO�G�s#Mg-��u�(Bz��	��˅ս����@m�2�@���p�@�g�ڤ����N�$`ս�#�G�V� �j��+�;ļvT�|��j�L�׶Z�8�&"��Q�tU6��X�������sRTY�QpBS6�^�$ ��]:��ן;� #���*�lO.��[��[�SE�HH���j3Q�7{�W�����*J�6籜�@ĉn�5����#LP��7��$FgGx�
[���&��Ö�f��R�t6jSK�����ci����!�ebdV;��o��_���m,h��4 ��@�Hk�; ���c��q\�~sy�r�£Tބr@��pƖi�B��3��,��b�Y�n��gXLj�z���W�~�Q���s���8�J�7U/��D~���tQo?g���kˁ5*�m��ĕ����0�2��!@ˀ���x�.���T��K�Y��*�A�+S�����N���9�^=%=@�%���2��J��������!�n���,�����x�.'���#hd�Pn�������:Ҥ�!'#�J����)P�I�����rׁF�"�r�a�_��=��jP�C�ͅf����^ ͧ�p����7ݐ=�,oi7�sD{dp����l�t��$p���f)�DA�P�oV7�_�|�Sˋ�YD��Li�q��b�z�Dl�i�I���Q���M�	gU;��O4���|*�Z4ﯤ���}Wv�Q���K��d��)�7�k}� ��Q��wq�Wg�)��*i���q�L�� �h� �I��M�1/�� ��_�<���G�(W0������ i?�҈�w]���\"���f@���T9�'����X�����,����*yJ��8*|�i�R����/1�G�ػ3�7�;%��`&u�v� )��;OB�#F vW�5��W����s>]�:�j\��]O\9�U�P9Ό�x��)K�RWB��§I��Uyf�cx�H������������� ���]�'�,�	v?�yP��Le�i����������<�p+� �IvI�BT�at�]�Wj�o���s;���3�dm��]	���캙�+:��QKv'���l�'�O�m����9���s�,l����?�S��z�5���\��>�&��z�b.)b�ۓ	���/����w6i�����S^ChZA.��d�)��E_�Iw�{Ĝ�:��7`j�e*_�9�a�I�As�s�FOb��ɤ�#q'z�X�N9 �g�z��z��_f�諱��ȡ~ƌ���{KC���+���b��=[��� ����RY��n?:�^���%�p?���X��D���]���Q`��L��ClҚ��6M����Qg�ρe��B�.);n$�>�>�Z`;��wb���,��].��i���ӷ�ZnC��x��Rǿ�U_�ܢ�$2��C� %�:���WXM$��p�!�Gp�ڛ���A��N�C���ז�,l�(�I�ælM�h����4-��N_��Hp��4�9�K/r�E�m���#�6����^"��,����4�ŬTGG���w[��u�*#p��^Y|�.����#�!��"~Ʉ��Q�\�`)�e!诒�8�4ycx�y��Ji��9�|z���� Z�Ms}�i.�L�+^Ac-��T��	M<毡�{��x$��"ǽ��D�6��6"�Md�L�ǥ�
)J��ٚ��7����t�[��a�fd�
�k5�G��t)��z.O�X�!+~��g���r�qٛ!*��7X��pi�?�s��	���3d��>�GKfX�nJC�2���B?!f���}k�:>�|� E���t�"�"�&�ɢ��*n�Պ���+�	���	�?�m:�a��e�e�}���.�61�b��@'h/qLˉ�"���y�S�I���JAc�O�P�������մg�U1y���[곐أլ�}ƨ*��?�ZK�9<�$>�tҴ��x ���q���M>�ڂA��(]&s0��n�҂e7���}��4����B���>��
3b�ECp6�©B�_���ҨF"a�&W;��~�@���X��m�y��)Uȅ,�"Q,N]Y%M�s@�\��:�ˮ~�}CA�~G���]���`Y�m9;חP���`�S�t���-|��Y�a��M��r�����|��BiD2״�^���l�w�������U��3����H(���,?�b� Ȣ��Rn}e���J��ݵ�ե������⵫Q�5���p��2�-
埠��9�ǹ�я����U�	�gWa�؛���U����Yd�	CX���Q�	�΍8�K�$g�Sz*FZ�M9>�uoU5��_�&yș�����A=���S�T_^riފ�W�8f] >��P���B�Ly����f�)������B`":��>�S>ҥ$���n2͵~&��⥷�LOiC61vS��+�@�������+�5�E}�Xu���ֹ���o�I�W�~�E�	ި_��|*ՁF�I�y���C���ٱ��q1ך;���/d>Pi�K����&:�,�2���S3�f���=����'�j�)�E\� �����J�q�\5vTv��Y�xՕ�P}��+�zY�?�D5�ݼ �[�
,q�C����r�h���V�l�8�:��iw� ���l}/r�R�È�&@�z�#�Ň6nt�QNS�}Q�_p#^K�G]��
��1�`ך��2S�YC��0�}�F�П�����u��)���6(6{��Ӫ0"m��9Xp�tm�>ˤ���\=����bC���۲�A�@�9��Aw ���}n�i������_6~�дv�O"�s�h�cB3��/��b�$>�EQ�_vV	g7�\О�"'���Ȅ�s�k.�")+���/%��������]n$k�;�L�i|�s�=�$ɂ#�+`1ԥA�D�z�@�*��tWѣ��S�D�sP]1�oӷ0���T�k>�R���^i3��5}�,lؘT`U��ǐ�&��w���~(�:[�}Jj";�����Ԍ"0��R�.�&@R��yHՉ�;����x�I3�F�}���Ps02-���J��" A}:Vɡ�C1k�꒠�ٶR{-�p^1��}œ ߛ���;�%
�#$+-�;���ފf�5yq�3�[�2�p���z`�ZV�="K�_K�j��D����6�4�+�<��\;�OXP:T����.��)��Y��;f_�0tƄ,`,�a��Ҙ[ĵ���E.�C�'���� �+F�v	1�M`z±0h5jos��^��klj�Y6����V` ���L<�n&���=]��-*�"h�¬w���0��.e�����cBۻ��q�Ӎ�zJ\����,�l{�q0�B�ˡ����Kc�Ϟ�a����;��U��A��h��Pۚ�|ᓎss ��g�a��k��QV觏��CQ9��K���X����ۉ2[����qel�~r幓de]-�9l���5��HP�.y��	�"cm���Y�n�7��E�Z3 mV��Z7�������\Iَ!G�[�)m��A��*SF��C=�i�S��zc�G�٥ϙ�(wf���$�6��H�m�QVt޾�E�,+�T־�h�����⤈�����d��n��Ǯa½���ķk8S�ɨ��)��%��`.��LE^�/r��&�G�����KE%
q(oP1fT��Q#V~�(���d��Y�`c�� �*9�r��҃x������?C7@0��[:�1S+�2��̻a�y��2��:�R)���hBK-�p��#�M~e��6��^SS�rW5�=����w�/]�s؈�lHeS�z��}�ju��N�dx�9��a|(��8�[�G�n�>>�"�$c��pp�~�(�ڨD��-�Ȉ}��q͋�)B)�p���2nZ���߹totVM.3 �p���c�0ZZ�$�BLf��5�����֗�����`��_}��>*΃����B�)���[]�Q��#L�~��~�O�{��۠�g��h��j->�WR��tG��|��eK�f�F���r��n\pc�����Z�!v7zn�U�����BU��� ��|�FѤ!S"u˕�՗����C@\�x�5Y��o5J�'2Eͬ��d$Ou���r�}����$�����W�7R�!��;57g��)�Y6��d{�
S/��O.����i3c��@���݃]Rщ`�D(��)���)�Y�ݞ E$�T�1ǅ��#,�j�,��.�eI2��ݴW|�c���Ġ�vC�і�U�Fo1�(͸�mߪlR<5h�$e�����C3x�e�,��e��"qZ�V�dx�e���Qz:H����q���s�2 7����.k����Ai�fȥ_��{�C�Z���A�7p:�BS)'�fo+�#�y����Q��;����b��;�9����y� 7�ˋ���"��=�ʿ����H�!�=�2�5�t��?+�+�fz��{6����d�Mf�|ˁ��=�
��l(��V/r�Y(���::2��?�B^���cP�=�!v���|2؝��\�)
3�>��0bU��6�QT�-��^u�7�L�Za�2e6I1x��5��t+�y���(�9P�2��UJa��j��u���b\\M�!m��k������]ϓkr�m��Ɣ޹�Z�G~�awJ���Y�l]Ә@��y��=�����6�ٗM3�o����0�H�X3��3{r��q��`����C<2G�%A�L�97�ז��iy@/o���
x)4�&������3	8d�T�	g�;b�������J�B��b��[h�H�����Y�6	a�$I;N���p��tnIᅙ8DH�vM��
�N�֊Lc�L
�)�"]}��o�dm��0��!�"���8'+Lp��S�Pd)��[ /����������'�|�?x�1��(vW�OE#p��E?6���Δ;��E3r �F�ko"�n��V���W�]�Fp�##vξ�1fv� ����=��)�����B꘹	P5���a���
�!��ӂ�T7���<��Ip�-�S�T�3��a��¬�UA��~�8�TB9+��`j�2�&�{�g�cwn��o7u��.�5��8���!��sﯦ٫�>'��N�T�m�
(+&����.�P7�L���/�C��{P F1�u�)�<��D�r���ɑA�l�aIyB]�#�3p��ݓO�tCe�ep�#&�߉nyX��RY���S*�؄��ffW�~�xB���#�kS)vV������e��5�M�54}�D�g��|JE�"/6	�޸O�D��g��a���(fifp���pL#� T%����8Y>q��Ad]�z!�(����m�N��vE�흔L�Ë⅄c�@��u�kX�����$��n'0�;龡n܈^ޣ�?.ǌ�_� �qFM���������d�I8LI��yKҘu��ĚX^b��r�p�~�@Cc��La���܊�v����iW���xr/�I�HԳ�l���k���-c0L���~b� �ΔWkC~�~�F6k���c�R>�U� ����R;?:i�xK-����Nh*��~_�e��G^����
-�Y,p��?��P:k���Qg���3s�#��J �����PAp�N:[C�*i�u����D���+0��F���9��J�b���]_��$f��D�lw�-���?�n��P��j�Mz�+^�����]��=���&�7x5�wG¯�O�XK�w/`-V1;X��kXR���1?Ŷ�.sc�<E��hk�Qb��G��/Y��֥�ltY��}$������\>7Ů�~6�*EA4�莢�(�˳%��Ǜ��zH���s٩B��U�yoN�f��>��C�G���8Y�3����o�����$j���R6����!ż��R���)���zx%��V������Q$դz���Y'5�4�0�����j�s�G�c]P��R��r%[i|���ʁO�$�1�8ʰD�ރ��<PR��0��l�DgΩ&�'A���yϸ�NA�wSL�Xc\Cn�tp����ь?zt��k,IwH���BO".�&9
�h��8�Jp���""L��n��%�pU(8R{֗��?���z`�?��juc���n�\aX�Q���~��Qޚ��\Lef0B�M�┯E4��KcJ9�"@�����=;S2�9�fP7N��*�X�E�ῦ]�2���/�5�┛&5���J.�a�c�(��,�<NM��<V�׊L���r5p6Q��)��ܞ_J��uBR�榃��2�^i�(�hʹ�=c{�q��xV�l��Zi�M��o	Gi��p�c��L��Rs֐�r�K���L��<��������`w#A ��Y�h�qԚ?w `��|�4����űu����u��n��P��W:sL8}�e��w�j���_�jd�NDdg5��o�]Ї� �`�-m�k�(]��Qc��w)��R���I}����a���� ���K�����~&��#�tGq��`[J=\s�$�`>=��e��=�>�x�x�R�<��DS�|��YhY�1C.[���M����{c&���J��"ES2	���� Ȟy.!�z0��J|V�ˆ�,��������C.�X��y�Ic�fM8���%v����.�+<�^��4����}���M$t��`���^������<H�r��i�J�#��p����f�P�V;f��������R9~Fx��-8�֡��(Sw�4-����ה"�EJ�y�[�M�bP���$AK�+Zt]B_U{��S�Qh>���)5��ivc�0�~n&�#pw�}�2ҡu.JM&���.�	�DtN��8.�SZ����6`��Ie���D���z�.�oD:.�����r������F6n�1;0ާ�<}IxѠ�G��K&+x�b|	$�k�����gl<?]�l6����5�E\Ee}iVvWle���Pj�9�T��rl��e4��Lm���ŕ����Wm��pG��MǪE{~L;v�a�TS�̳�JF�?�s����D��K�C���.��;\M+���Z.�x��Q��Ǎ�Q��U�xˑ"��T�W�",�C����w&��8Z�O���"�*�⮍aAS��v:Rs�="U�a��1���J��G��-O&W�ĳ�@�b��2[�J�^K����r�d/&6�ta�?�D�����|�aB1pA^LV�\������Tȵ�� ��T
sh�S[D��X�Ȳ�P]�W�M��ed_��j�`��˲P��3S�̻�N�;�E�>�Ռ0v�Mױ@������7�R>��s��fbr�u�)����74����c!��y����/
]�����\_S;4k�ۜM�e���N��\��iU��cCk��74_�`�9��;���՘��S�
s��c�*x�K6�ȗ2F��J�ˁ�B4S�9��������z	��Cm��ˍ�!7m;mY���>L�m�k���.�C��*-��af��|� p����ŋ�e�Xb�X�W:cb(H�ѭ�Ty04�`�Lw{�x�D�5`��\{O�ّ�]~L��z�R����(��p����`18�Z0�S�%Z�����Hx�J���O���(:�`MDŪY���Y*�W�)���O�N�%e��ۋ��W�ֵ	L�ڋ���Ib�"� M�wOx��d$�Ǐf:��[�[�+p�T�r�T�ޛe�Hf._uO��i�>���區�r0	��W��1���F�]ǂ�$4���m�(�Gvݯe�ۻN���$�CBXv-	��p@+���|�O��Q9N��g�8�t��Y{��>�ro��������"L<���ݙ�����u��>��_c��'S�6�B�f�j��X����bb���=�R�WT�k>�^��p~9����>�79�D��΀���փ�/L���|!ؔeB�ܶqxЌ/�֩��`����jB:X�2�~��U�"!h����9�߃�;�_�D�oF���L����EK&������k�~����,�\Ẇ�$�J���V~����p����l�G?�{��v�"igyV+��#�B{ ;�8��Ung�*]�4��T��pMR�Zq�������$����Y�m����ot�V�9�Q�7����v��/�6���{���AJ����X�����C�_�6�#4�Ǽ��ixktY�t��V�u�C�_l75��e�
�x��/V~nC$���~:15s�H�����5��?KqH,q6츲Z���hT�����0B=��~l~"��z��O��w"��������yKL�D2��N�aX~��#��_6ʸEѬHy�)����(+�j3�,���<�'F9V����� ^Q�H�J��gQRR'(;�	\�PU�mNÍ�h�̴ź,�ȓ��B��7v�i�@t�?�/���������n,b�����L,�ì5?����e�!����s �����򧋺��{wr9���
���Oe�Ͽ��q7l��?t��hc� �	���kL��̠1?�^F�t�bAwI�������㸝F@q�B�$N�u�����k�Wӧ�c������%ce�Hl�n�(�Ih��g��&T͔-����J���(��Q�#8M@wVk�
~t��3#|��j)�{T{�7��g, Y�d
S|���+k�^��W��qT2�Q���x�m�ȷ�`�rF�7E;{}���`:�J�\ж��j�pv`u80�"2u`���w��*�6�b/*?R8��/���(�}#�V��Su4T?����4�~M�y[�s��Y���٤+�_�J�-3�a�m�j��"�<RHzv6�,I�A24��#4����|���k/lk��S�3����I�	O�a�#R�!x3�*Ɖ��(2$��rI��T�1/0�� ��|����N�� L�u��J���w��:��ݒf�zq�OtFQԪ:���MκO�I+l�dN��S��T��.��8�+R��}w3��_L�<nb��+]���$���W	 [��'���)�\�嬎�ԅ��<3Q���QWJ�ȏ�g��I%P���� 0�*3Z��=�2ràd}�Av���G��`ǫ��?O��Dw<'�	�6\��-}����|(?[��;�  �:��S�d-�3Q�k�ccεJ�j��JWp�����I��!ؠ�Q��ua�"3�D�^1�����7��|����q-L�����%JQ�or�NΔg34~�pO�	�߹~�����ց�8��ҩfUuP�J
��ϥ���_��0`��
z�C��t�=I�q�j<��b�by���軦S`0KjcNj����8@1N�����p������pEr�A�s��6�Q_������'��;��Wh��ij��4�/�h��ᕮ
�ۺ'lRy�J�L�nmc�B9�Z�q��֩Q-4�zR�!s�P� o�u%�&J���{�������,Ѻ �$�y ��m�������w%x�4C��F��C��m������W1��p6!�Pf�V^d�]*t^����W�-�!6�2�Ǔu�k�7�� t�=�:{㧔�����@��.��h��T/�A��7����\�1���߯`�����=���k�����m����Dy�>�[0o^ om|�r��*�{�ctL�r���mW�)��>n�3e{��Bxޡ�,�p�;�2��e~4+a �$~T漩�
�����H��1��E�Zy*\�?�|<��
o�Z}�^:ʐ��	z5�т=bkVj�sO�`V|P�(@>�%LNBh��o��=h	m�C�3f��pw�!P�+_c���4�o�Y$N8���� s���r���_�٫��Qu{��E3��`�D��0k��Q���h#��;��O�/�gV�e�s�iA�#u�g�Ķ�i��m*nH�9������c��	Xp�;ӒB�,�4j �|�uĂ���~2V�[&�H-�~u``���B�����W`FS�lY�4v��/x��i����j�g ��q�l��"i��k��0s=Y� �2�< ���R'�ݙs���FH �k��Ya��J���{�yo�JKtk�%=N�H�+�~�\�͜�B���1-�Rw;t���Z��gb�7��wy��vc�<&ގPs���ⶺ��.�����汬�(�͂��dR����Ids�N�6Ȫ	�AL��Ut?������	\���C�w��`y����զ�t>��ì������{a���8�{~�'�H�����]�ȿ���Ƣ�Cw�1r���o4�YЄ�zVnq�7��>Uz�H_�=��k����� �[qb��7�vQ{��.u�G0�B�J��zmU#���D�hڋ?ȷg�46�{��E�@�u���@O�&_�v����X!+"��m�:�R�לEKF)ꖵV�uQ��U@uj�a���g�5(>�"%���z�?qكu��e�b$�$�uK�84,��\
e �Wk7����n �޽��V�N��i���
�*�AX�4���#��	���-^$���+O���j�Y�6�'��)�1iع��m&a�F��)�@TTܛ\X;ou��Ock�Xr7@�������0Jx�0����L{D�q�E]6&�z����m3�����˫�EuThJ��!(*�7ޑK�}4��]�nF�[�9$�9o���̭�i)J�w˩��{�T�1��h�f��{̍&?��c�-��ñ@�;O�H$��y-z:��3�I!Ң�j�I�,����c��Ql!+Zx�#����C��eh}<��nL�ύ���-�?͢�DH�f佶��oC}f'�RA�d�M�j7z���i��I�W�B1\�#�h�����RM���"uމ>T�U)����M��&g�XU�0�d��_*W:�<���#iGA�c�@Q�􌊏&�q���_7����	?���vѠE��/)��'E�q��!��Z�)�$�0\�
TXoCP�̚c$v���G�ʩh�F ����1�����vmg%�4ɧ�~J�����&�k��h�f��'^�EiW��v�_�M���љ?!˄����MW�]��ï�eB��4��F�)>,S�O�G�����n$Ǌ�����a_�&�::�f��@Aq��b�R������I;��ʄ�O��N�g�z��̱�9�7}a����0I�s���W8S��m�U��c+��,��X{��㚟�A��� �]�*�K����yۂ.�=� Y��=My�O�t���m�R�����F�7w�g,B3�?Ja���ϧ7/���'���$ƌc���a��k�/���8fR�8ya=>l����3φ�X���a���5sˮ�f�n+Ge}��U��:�%�pm?��*~�%~�O�g1�h/ߔ�7n�yЯ$�Ĝ�F���?�c���S�2��&L�����]z��鋅�<��H����3�Pgz]�(2�`p����h����m%��<�R%���Q�y�f�t<���7k�w<��L���9��	0�D��|0'V S�d�MBz��_ad�;2���~b* ^��<��C���P����M�AR@OX��d�t���S�IL� ׾��;&f�0��4�w��u������-�$���9�_�ު��ʍ|Ay�Ρ&��N�a�1_�Z��l i
5�
:�v:��Q�Q�P)�p�F���K�d��y�3�5v^�Iy&�:��ʽ�E'��t�E)���B�8�X�ʔ���ʹ���Q�#�C�|>����(n�Oi��bl*�RK-9B�(���Wb�\ph9���~���:��O��W��;��!�9,�z |���<��lfL�}�b��F�sG#q��M�Yx��D��� Vl�ZAc���VzL�gL'9�o�E��"��zI}����V_��̀m���Kk��bG�m�aX� S�������&8��ݩ��M���=�rDv�<�nl��{#!Ν�
��oJ;�l��o�Ef�ɒ��0�~�����%���W�9d^���N#��*�*=������z]w�$ӦJ(N��`���jI?��.3X:�����c��/2@���̩�[�;�Zo�,��*f�nK�v(C��CKǏJ����îJ [ k ]"�"��Q����0K�Y��0�c������I`��6�S����� ���A�旑�9��V��X��?�pk�Al62�:���!s*��E�ʬM����-wU����C���a��Z+�<�IJ��"J�J��#���&f��.��w$���wӴ�p�Gѻ�S�Q?l)�Z�LK�}$�7����7����Y[���@����M[
����.]^$Z5 ��k�##7p�K��F8x=�<�j߼mѫ<{�[�x��<����,@�����n�g�L��C�}ē�n\���e}5m9�]e�~E��? �s�S��x�kB�<�|���B�=���zH�%���Nf	�si��^m͖.��v��K��RkG��E���8:T��j��ݱ��^1J�����q��}�3��IN�h�YPFB��R�9�����x��t��Ӵ��ϱqS=�5l�?,5f�~` ����,��a��^]�����ɐ���7�G��x6����J�n��*�h����G`�xr]a(���%�L��Ϧ��w�\�nɔ���C���/)�q���mt�UЀ�<�A�e#I�_�l�5K>�.�.#lev3��<�[BC�-6�y��[&n&T�����ﳠl��^��ᦝ��cWW,�t�*�#���'��c�_j\���u�g:�1�-�L���yǄ���	>xu������ط���N�r���6I��&����,]��Ȣ�;!Y:��dyS��x�v�v�����î�tc�~�Q^E�X�rDu�����Ch�-W�������.p��N�yl�t7*ж�?�r��o�5 �:ugn��1em8y�GB�&�J��$���E�N�^:l�`���*i0y#ah!sm��B6H�-�|��/�T7�VOTl�+����.:hf��6�!4���z�Ե��U�nw�#����`%.���_'��R�����r�'	<"
aś���T��ߛ�y�ω8�� ɗ���6� ���J�F���kz?�5�ҽ��oMU˽Z�|����a9�'���q
�E£���)'SN�9�7�R9g��a^�<p�@(�����
��F�/O�%�}za�j�v-Jm�ƅ���gб����n����T��tkhlW:D����Y�M@���H��v�?QW�D������O��P]yT\B@b���w�� ء�[I�t��C�k��m�b0��%�����$ �H�☐/b�]�O,�~�Y��ǫ�A~�?%���v{�g�W�Kc�?���b�uw.�)�	�����~$d�1f���OD���H�*�ǾcJPͺ��-�uق+�)B�X�Ȭ$�u��i�Y9s��猦A0gQ}Q�I:�v��X(FW��~�z��u�A7C��R�m�D�u�xJi(�RK�H�I9zĸߧ�W���рW�,Gғ8�[�(�.���羽�h3S�%a�F���b'�
,O	-�>\�o�L4ȭ��������y��1$��yi�}�����T���`Yf|�����w7�:؇�.V8@�ı$/�U-)�'iZ�8:Ռ���2�G
xl��hn�%��r$N��P;���������IA���2��ANm,�vK�c+�l����R>���*���
R��(�kY�/'���8�A;�"q����M��斏z�8�����(�Y���	8-V�=��fgR$yXo�f{�H�ߎc��&��6�:�{퓉�r
�j�ʒsx3�xN��j��$vV�-5F�(,�h9Ї��6^�*��!a��O��^of��<��}�<�F�
�D��Y,���#�q�czo�8,��+��X*�d��NJ�zZj�3ᮚ��]��д�ӤS3Y�3�cQz\���-��\��3aQd�]7d����ۦl6x��w��y^ elEJ��ݲG��7b�>�����q�bw�r\;Ԓ؃�Zj�iy'���y<'M�i\\ 4�=��a�D���x���� �%4�"�x�D�n��@,_T�E�"j�����>6u��Mbxj~°�r��<5V�9��h�jT�U`��M����JYh���sI�m	`C���b*��]h�7�73�=+��RS���-ψR//|�4�r��z%gy$�f��"2û\a�r�b�'#��(�3��*.N%b!�sx10�d�>'�PZ�b[��oh9�Z�}Vv订<��NG2��n���/�dn�@_��E$�QmǄ;t�v�������l�}bCf8+~�!����N�,���4�D(7�����/�D�¶���R �al/���N&l/'6`ua$�*�K-#:bdE�ub���5�ӗ��<ڮ2�$�Rw�3Bd���u�6C4񢠽#uњ[ҵ<QS�'df�!�\�I�4W��a7V���1˹]_�� ��ߌ��I4 �w��7KFu2�S�p��L�+�߾f��xW�6U�0��4W���҆G��#E8y	�F\UJ+N^@bB��1�atl$�����w�J�N�!$gd]3س��p�ȍ�S�8���]~㋲�zV�Tu�"ȩ(�>�>��&�F��}_n�Hԡz�t�~m:�����n��#��T9�Њ�)O�|�/@�����#��@��dd�� F����)G�-�4�j4�^b ���_��?o�  cG�[w��
o;Л����A�q@BÓ�ٽR�!4���]�����EĠ[ �Ҧ��Þ��/�����$X89q��&қH	l���ؠ
Q_�6����:B�9b^��2�KH���R'}Ґ��I'�﷣R��o��F�������d<�*��Rmηd8��:�ߝW;��,�Wԏ��j�O��7�~I�;��'�	�>}&�9}��'$���=)���K����0R��� ��6��B��n�) �=������!��3�"���qr���@V���'=&a�}� ]�I�X�*ت�����"5�ݐf�|����Y�L�j�WE����1uB'��i~���Ia�*�CNN��Q�;7ʹ��xG�����N��8v�]��$!x����A�}�UVMkȩ�SQW�٣��-[:� {��ىots�7#�A��{F���U�=$���U�+{}..���.:���X�1�;x���[Z8���:#5�9�Hy]Z�c.���T�!'VS�����Iw�^�.l��j�T�L0U���$�)h��@�D���8��û����/#�ީl9x�Â��I��s��ظ <ݹ������[�� �s�H��x�Dݏ:�.w,�R�M��I���n�'��=K���%e�z픍�mΊWphh��q˟D�%���b:�8�57K۠��
N y����}�J��2��	�@^[��:oW�;`�.,<�qa�z�/l�ui?���g�y��B`�j��Rd��f���!k��ZT��	+~���xm"r�� ��iRN��<*������Z�o��8֟7Ť�R"�A�TX/�Me������(P9�*х�k=k:�}Os�O�5Ryj��8-;���αڞ����I$�AF�I�i;�"���Xp'��Wc��Bm����x��A�`.WO�c�N$_�x�V��ئ&��>?���,W0�i�N�jĚ�)d���v�e	��������q�#�+����9�ks��^w��8�U�D����w�5���Jq5{�]����υX�%��V�n{�d7M��aL�d��A������&ԃ�$oU�2��7	;C�|��g*H��l���d�*�y�`��>H�ɰT/�{!�my6��M��ؘtǨ�Է7��Q�{M���Z�\��:�CN���︵�!�Oiғ�Bڽ�.B����l`M�V���a�~i+OU�f�%`0D%y���-ĕ��|�S���n'�Od}Т5�!��V::!�;nW�_'���e�
�k��$���1O�ʰr�g��yHg�!e��,����y�5�P��A�\���=jN��<�$2�ʊS�:�|l��(��"i`���J�OUg���P��<Yܴ�6��I���P���Vx��-1{}�e�n�B���CCl��"�N�VO�:�k��� J�G�9D\i�N�)%W�=%׋��4O/���I��lo�^�1�-)U�a㐟,޲F����E�/�|�����?w�;�� �����R�S
��RCK
�}�l�Z>�d��ӣ}<�QJ�Sw��Ծ�rRr&%������t���K�� ���� ��Ф!���.���
m���N����n��v&�H��O�1]U���.m3��9�����6�B�=6 �N��#��n�qX:QB��	ҺuxF�̨��h�
���a�о�Wk���z�Eq
ܰ�.�7�@6�pw��2]iA'��b�����(+v����,Y:gի�w��M'���7x�^z끅Wց;j3�p�Ж�`_@Nk�(���\Jn
�ZՂ1��/�"pB"�;c���'8�K��f��T�*7_'���}6��F�Ct�L$ ~�nP[p(srӎ� �ľO�D�D�}��'���� .�Ԙ9�rZ\��ʭ�yQG�,��X��;�M�������!<�3U���qQ�:.�9�'fb`�m!M���m��ڑ~i�X�D���)8�S�4��p�1ְT�Y�pj�+�X43�6�ZA8)�������`�&�V�yձ�l��ųc)m���Ϳ=�=�J�Z=��4�됤���lP_��k���Uo�m�P���b�>;,���2`O��������Z�	g����6l�nw�qZ))9��
�\��l}��ۢ���o��G���7�K�,uiX������K�&B�i-y���kA@l6���JX����vg�7&�S���j@�j�g�4.�B�=�h�����gu�s��۠�%?ވ�����72Ir�/�-..���>84�]���]��3*��]+G��#Ptg�d���Ǽ_5��p۲�1�MW3���˩�=s�ZP�<H�s�r"7�Zh�]#Փ-�;�N)�N���c�x�|~[c�\���W��C�p��e�;~T[�����˩���[��}$���V]3��)e��Z���^(9�Ť)֗2�?��B�����H�U�R����m���HOϱYK���=BD��QD��ke���~?2��O�*@2IrlU�A�DcY��A����>�z����TL�@tʭ�k�3B�uY��}��ǒ�Y���S�&�pg����e�N���&�9&
"S9ƕףI��VJ�v^��}V�>62�&�yXKU\2�����୵�'����p��\	��i7���W����i���l��դAP�(�6����\�7;���yÝ�k�B���)�I����w�c,� ��Q��y��P[����K�`Y��N��-0�t�G����[�i;�0���V��
�DI�*�ͥI
�=�����a�c�z>;�|�K򱃩�������x�����Cx���_!��"��3T��ee��[b�~����ƜȤ[���������� ��*��D-���m�hN�8YO�{-AU�E�l����^/�gg��8kR�;�w��k��z���s.���E<���C=���O�C}�Q�P�٘�a�/vO�>�W��
���K$�^$�B���~�1�]u�y2R��R�/��M�2�����'��� ~@�����*�yR�È�Sel�[K��ij�|	�06�"���ȢǴ5D�C3�oD&��>_/��b6�z��@(�luґ�񊤧*JtU�~��S�z8E���A�7�:���[aT�8~T��k;�s�P��dZ��(�+i�X����<��|�!̄�r�+�W��:�7�A6������g�u��v�tx��}(v	M�x��5���o�1�)Z��8S.Q J�e����_��F�Ϥ��~��4a�ؗ��2�ظ#�;�����E��.�B�h;���,M�Y����;j��_D��	�#��ECJd��?Kh!a�o��8�ʪ�Z
�0{�p~��/�0'Tb6�@e7?�fF���h;��tۦ��-��u��ds	�'��.��|ʅA�O����~`e�1�L�+���3�HȎRJ�}�Of�I�(� �N�a-9������2�b2Ꟛ8��!>�|q�M���Hm�\�L0���|�3{���O��8jM��J��I�}�Zq�q�=
�0g�ȫ��-dZB�����~a��l�"� ���*�,�Q��Oc�i�\$���]��)�55#Ǫf� ����hrOA�`�}��*��M2v洟�|a�,.n��l���lO�����{*h#�z����}�«���n�K�������8��`tb3ph��
���}�b��&.)q���]��Q0S�j�ńYX�����̴�L.���_��7=�o�kc�9��1C�A�YwG+�e�__�^�2~�I��/�ۖ8[��T��(3P��s%g�Ĉ��?0�f��;VGd;53y6v�w���4��߇y%jb�t�-����2��6�>|7uν�v�ݐKG�!Ӊ�DKu,o�"��ֳc���b"�Q}�&�PbQ1�/�<�b�n�E�`!ĵ�g��J0�B!�9\�:�7#-�[�����W�ټ!w����q����n���l�����/BeU �,Biw#a�2Ρ���w�*�4�����i�r(jqz�Jl�����ԝq�� �U<��!�V��h�MK�j�=��
�����Ik�)�Uq�[ dx�}c��k��T�j�/L��o�!�%��K̍/��|��/پ��=�N�Vw�Oߙ���@I~z�k��Fy>ͱ��]����8�U|DN�n�h��������Ϗ7�I�v:�h�F����K'��9����*X0�תn<ƣ�'�g�&���.�kl��3�&�`��(%��eȵo���'�ݳ���?�!�!�&?B��c�����z��d�.�>���h]����
���K��x]-���q�2�So$���9��Z�B���L$$�bVE������v��s�%&T�����G� ���t����)S���uC�t�4�,�&/�ma��3��L�l&�����;��Ds� M6�*���L���9h�p�6G�Ub��>��r�t�o���PJ���r&3�0���l�Vp�_�d#��~~�ub3d~1No-E�^*���=���%H ����ǜ��#�?��ᑜ������0rUش�/�K�Fk�'H�b$���0�N{�(9�꺈-Kq�gԲ��ATz��5G� �@W��w"�`嵗��<[�ŵ�
N{]t�u&�K�0�7z���Ꙑ��3��"D;o;u\zDt:�3�F�n�##�������+�[���ļP��A|u:���P�Ņ˷�9�-V���I�O�&.]5uR[n�����Mo>�� 7�Ifj������U�K����π�͍�M�]٘zPW�i�R59��'_*z	O��A������tN�v܄e{B�۔�2a�&��6��̓�����x{�{�{��@�@�+�;� %���Jͼ�1FP���,���V�:7��%���hln��wo��&ѿ�r���It�-�aaO%��/����:x�X5��/��/��WTЏd˩�N�kR{��T����z���r���$����Lؓ��J��ߍ�Y�1��ȹ�v�c�� m��|<"p�p�f�{?ɣ�ak��#y2Υ��҈�|�#3z �k�x��tL�����G�=�l"�5��"�O�#_��n��S1�~R�f�n�sj���9�LC��r�⒧�sI����!W�x����-B�0��)?U�$�h��������c	OFj�{V�.�_�O��V�;A�}���ɶ�|��j4��p��,c}풼�����.��@��{���t�iTu�m�<4�W�]�0���+𱆧�?��ۇ�����1����@XP�'��yp����B)R��g���S+ko����-p�Tk���l:>A5v�f�<�ůo\���ht�J�^��aj�Q�bɡ�=���T��OU,e�T�`��z/���C�~hN6���$��Ե�|�N�M�r�������	�=$T�W[��	m�cj��)}��~�a��CV�dA����g��P~f2\_eq��B1`z+#v� ��Z�1��� �&Gn�����J1a�"p&�澕�di�[�>�sX�n,8�P�0�"���K�j�9�ʔ�~��-��w�{����c�����f��R҈x�7{�X_��{E�n?j�����<�zN7������΃��<2Ѯ�gI�,Y*>d��&���Ʈk�qnո�'��� B�֊�����;���
�tԨ����v?1���[�K�_��N���w�4\�Ķ�>D�;ŉ����}T2|)�{(�!�""��R�w���.+�^-��m�oB�(֑ീ�2�ky��W���X��Xx��=�b���B�s�=8'(wBm�t`4��yx�N�n�Ǭ��c�_�I�m��=�w��4ʩ��p�o���0�p�]`i�kk Z��>A�����v4;*��d��"$@�-���X�F5Wv-s�	�ZY� ��w]bE'���`�M�0�V$m�h�,�6��:���d)1�ü���J/�|����-x(+0&�����f�����T�NQ������l|���&��}ϴ(p/
�Z
�oƞH�������ttTf ���m�)�0���wO���5O��F�h�U7�͗fJ�`���š����
��1��5�L��I�����0X[M4	|�u�z3F3!�B|C`h��(S������9t<��~c
%6��Q/�����UX���.�
Ko�Ũ�7�O��y��i�vM�5e���R1w���rt��.�.yݐ��-�u �V�o�}�~(���4���蠖��"
2l�ⶖ�٨�_���)H��n�i�Ѓ�����9x��\����kIhid�d�u��x���Ϣ�;�����J�A]�aͳ�'hm�5�[ٗ#��\�=�9�g�:�]x����F�Z��Ñp��Ss���9
N�RK��C��]����
��Ľ�EZ�5i�
,H��'�s�VϤQ��)�N䇋X}�ʎ����c�Ѹ<o�"�<����'#�04S�)N�(��*�2��,�$��i��A��"7�9C�|�Զ�ـ4e��8�0�'я�2��B<�@�M$�BY��u����2'�N�V=8: b(�0�3k�{C���P��4{���}/Y�;'Bp��>E�ڷC����%|�n;�9�u+ٯl��c��40���+�H.=+�g�����33p�9��+���.̈́�";��Rr{�Z=P#6��\�ա�.�M����O�Z+�R_�!.y�_�kC��V���*�ˊ^@��t+�Y��	��Nvü�=З������\�+sf������K��̐������O���:���8t�l62H,({i�YRZu���"�8���⁓�K��9���:���������r>�'���v��Zb�=ۧ�[��4LL�������,&	n�{#��%Zg�A��<�M�	x��QL`~{QR��(h�o��g�T�W����RW)��abK�E����Џ����''��S�0F��1������j�3R��95;��_w�$� ��ϫ��|�.��&�Yg��Ft��EB�����Nt)GE�IF����*Noݷ��j5�����S�[{�S'i����<�:R�Iy��<��$�r x�0+A`��>�Q%��y���qI�Q��/����!�VQi>dm~�p,�L��z�[����KL��"�S�iK���?�PUU>�e3��LZ�)JEd^��=ݸ�'����&�f��P�r�{��Fw�}�8h����v�D�����UH锚*�؜u�dl����B������+�ފ�@$�ۧ�ܿ�0,'��	E��̓_P�5\*���C[�j<r�d����@[G�5hE	
�Wp�-��*�(�p1��j�tg�6P���!$��B�ѻ݂���h��z�x��a� 0w�\�8C�
Z�k�O��l�W�������T_=�^V;U���-��ʒ�]�n�-&2UD�]�vZ���&Q�v�^�KW�S��N�e/����@��'Dn�.>�1�9A�^˒�٣�S<��pN���@��l�i&g���"��J>\��&�^�	���=�!���!yM�VD�ɍY��w�_Ґ��t�ՁI@�L��۲�o_����mJ\꼏�p(J�6zn��4x\r��uJ<�"��d^P0�~9h��!�N_���,kY^)*t�~4�����?�Y����=�p:f��Tds�����S
R�f0�{���Nɲ�z�w�R��T��$yPu�ZK�I�"o�~��纡x�����1o�Q}�Pe�o4H��?B
H�+���!�n��ek������I�e Si�|�i~u�(h��*��IGU�o��]fE�1,�
���#b�\��<�כ�j�3���Px-��0Z���,�u;��<����@�DJ�n/�7���S%��ݐ5Q9��̄%L9��:2D��Săt"�4,92��b�1�8�v��4ݴ/�����׮g�tn�0�Б��>��daN��U�nRj�l}>;"{�9<��锦���Idb��iH$,��GZ:��tr+�U�|��X�`��>n�H�i����i,1��%4�g��@���\�m
�����
ClR�`��u����FTl�ۙC�?</���e��r^Y.�cy��O�H�]U����[�oA'C�P�:�%�%a�~&�h���?r�;�YN5f����L�v�F�S-<�WAnc����$�eq�f��i>`E�q��1���J���
[B��O�ԭ�} �>�)�	��d^ �L������K���e�Z_�o=��/�h�a�x��}����_��p�yrNN���ۭml
"鲗<l+�9�\�ޮE�Y�9��8idx�)���e<pDo�S�CzM�S����O�d�͘�Maj��[��qWTq� ��-Д+w[�9��E�ɶd�����e�bB;���)S�x�6H����4�*Z��Z5����{���s*�v���B��3�j��82�0�F�\���>&��#vQj�b��EǠ��?͐ ?����܋N#�j[	H�k�>�Ꭾ�0�I��N`�̃'(��( ��΂r�D�4�p���2>�
�N�;���M���%���#ȅR����Z�<P����D�#�0����ǁZ)��f��{�	�MT���+y�p�4=��U�]��z�i�`������A�7���F�8D���з�v��g���3�N�6��9��jU�H=��Ch2�Ża��5q�{��ub�N	��s�1�����Pq8mo�Ã`���w�\�0p'o)����8�v��2*<M���&pAqDM��5!ȣ�ئr��1��xc�D��9��k`��<�h���=���B}�Z~Z�L�~�/�����R��ȼ ���(��e�b.FE�$d�� J����F��
��1�$��qV��*�&x�C��8���خ�U��F"�_T�iԊ��imP�F`����\�YE�,a�m��&s!�ߔ���vs&9_��*���X��%,�v��-��Y52i7�6ާ+ Z�<R):������%�+�,���i4�XZ���R�]�v�@bJ��"���P��=G��%C��7������E+tNdF�S<2I�E���0��6��X�CYI[~i8���	���Q����oiEWA^��`cv��Y@�WV�v�ԝ������/�$Ǿ�1���1"���r��:�1���BҀž���c֘i(��u�9%��@@9ܖe�:�|�V�
���H�mO��3K��ڧ9N�g����u�@�7��QS˛�u���y4GI޷'��E���A[e�ハX��p�~4wW�؞�	e�/ml��k6Pd��ʱV�|(r�g����g'���A���!	�a�礨����/�ʃ�g�����P�E��}�n5���w���n��㢅��EOeZi/�݁!PN�
�Cg�-�B�Oy�L��]���˭}YK�ӈ�M��^� U���I:�2����8�789�s�D�x��R�Y�K�7�
[��C����]f��p��1��m�t�E5F)���S� ���E����k8�`R�^�Wk��Q%et<Ybu�M*4㒩g?�5B��1Wdf �3 VB7g'-Na�'��t�O�%�ՎĄ�3�y� 'b��|���|���s��@��+>�L�Y�*`�;�#hc���n��
!��k���q?���KlŃ�R3�@N�՝&�N�i�YE?ؿ9�������ݿn'��S/{Y�|�h���{���{ސ�Wt��P�	�լ��+��g��|ff�S{"����ԠS�Q�%��M�T�n?�.C�,�&��I��ar�bT�t��$�2�g�������Jue���|Q��n���C�W��k�h������D��N�C=��@H� ,���s���&}�|�~��ku�~���#/.v�U��]{d���x'T��z2X�M�;�O����+�����4 �����GI�ſ᏾����p ��\��#�B�GU��m�te�<���o�J�����`�$�)�>��6��rS2t��w0k@$�*Vm5���B�zu]���z'�3����d��� ������bg����`b�[V�2L��]ɝ���
F��S��/:����$X8�q�l�/��$ڢW5%P܆Kz{���B�2r�I1�e�����ݪ��h��Ο�T�����0�}�?f8� bI�ma�|�2R/bm�j'���3��gl��H�قss��K6���d��R_��B5��:�d`�y��f�̰Ƹ,qg���?�L�2C���v�=;n��Ewɇ��=�kż��7���.'��	��E����gK-P6�E�A9�Ű���~�9�$��kg�{��y��ED�;�tx�Q��T�?�Od�.��������];6�uIEd�q�m��x����'xsܧ�:�N��?w!���)�q�z��F�.`�
���W�}ɘ�(�vW�:g���r�Ҽ�<Yl����z4h�p�-b���&F[�[
�z���J:#m��ZPc��}�?]��W�lD�/BEZ�ehE�G���뛝8�����Aj��8�O+���k<�����U�#LZ-���sώR�G��F&����ϻ�����A�`�Y/o��3у��mY��I7+V�����h�7Y���c$����8���61q�����I�|8�2�|�A7�ײQe�'Ht�����h�L�i�����2��?��邇 1��� ��{�Љ)��SY���?\�@�sW�S5�I�.�kyt o��B�_w�W.���ڃ����ОcQ�CJ���5w[�_x��yHm��U\z��&����K=�p�ux��~� ��Xά�1���^lWll�(�ؼLp�"��UI�{��l@_F��r�I��d�`��V�\U��.}z�/�梇���92������q���S�V�r��ur�6'>��%-��N�ɼ����C�nt��_1�<A�֞;_l��#z�q�Ex�;��i�0����&O \�;�Q̋w҅D�W)U����.��2��D^]:W�=�a2n��6���(s�y���-z��m�H(��F!��L[,^�.cL��ȐW�i�z�Ä�hsx�k,��{�=��n��Q=�5��\q�T��Ɗۘ&�7kH7��'-B낝��m=�E
���*7kq���k軎������Pح���7�X�3k�
(R��!���:��*��O������M@�jϗ��cۈ:�ZgL/
wO:���)3sq�>K������|k]e@GObM�K�pG���o4�pUg��G�I��~��r9o����U�o���>D����:ǥN��I5��TiS��I��B� 9����� ��n�:E�mq�<{�R�5awQ# �f�gþ�o��}tQ�N��A��Jx�G(�"F�'�M#�O�]�q��uY���?������uC��I�����P�-�|s�w�nA�:�E�����.����!��h��Kr��b-\��m��'�D��:Rx�����IP-��v�\?!*��=Xo�	ަ X��!\�yH�&9�s����rBp������������=�y ��Ԟ(��0n�l�R.X�;8La�ӹ��2B~���w�ڧ�#l�����DրTpm� ��!7iʵ����� �O�L�N|Q���r��gZ�' �z�&kP��S�`=��p%��Os-�f.cjs�h1�L/�V�D�_��$e�����_ו"����N�:G����Z���h���*ˡgX�,�\eO��P� �{:�іwb�6u)4�>%F�+>N|r6��_
����;-��"��g�t �#�?%�\�`R#��RP�O�O?>��|K���Cb�Y@�q;�C��
ky
o^��!0&N")��h�|����tW_�HǤb�#����ɞ���ҳU���Q�B�ƨS��&�_Hi���Ξ��H�*���iL��fhd�ơ�t��~��v��)��Tq������,���s�wH���i$�:ޱ]����\�#oH���|�GW��X����ґ���a�+�Xvv8���}��U@����i��n�\�Y0T�+I�ٹ�HSE��R.�yiц'�c<�m5E!@(փ�E�.s�������%%.��Zٯd���G��=f�����&��.�˟iq�� �3w�ƨ����5����]5��4��'gG���j�)�U���M�=�I����K6���9����.�v�⌉����2�Ǌ����An{)2�hD�� y՗w��w��g��c��6-�m�o�P�4�9RW~��F�4�ξ�:��y�Wa'����ҭQ$c��U���%����mn-�n�T3D�"G}yF[vs����i�ui[�(�4l@0M~�ېV똓�7|� M�Y���XV�v�9 W��s�0:fRM?�%�?�BS�֞�*���ȵ���d�|�9�R��Mt+��_t������(j�⴯�W��;��=�pp+3&�t�0�l���p�W�V��5����u�0�R�r���-ˈy�"�C]�����_��:ʖ�I�C��4k�U��8���,^�`�}�mU�aH������..y wݧkl㤭g�����#e���ߛ��"KF����{>���_�o1��aC�%Lؖ�9�����&���JN�r����	0эz ��
1A��M��2��ݿ���� ��6��uL�O��t� �(;Ppb�Iښl�l.�_�uU��,�5)�!��V���@����`7�>l�����r��4!��x�H�[������^B�+�{��p���m�G�z/UKKn��Ӕ���]`�eF(lCt"~���(&��
Nc��^f�p��U�`��c�v)J����Z}�"�^����6%{K�V��{�	�ժ��~�^Ǵ�����4FT�6�lDKS��ۜC^=���V8�UO��d�U�� ���w�n�[�W)A�J�V�����+�%½��˛(m�Lu� u��_851y$?�Ff̓7�+�n��I��Vh�+��w�e|�>2%�p��M�~l��r̷n�p�N-ƤW�=��=�x;�_�\y#�"*E��ڸ�-P$yOuCh�˾�;��ٻ	r�Ld���y�w�`��bJǌA)�kp>���T�s�"?6J����P~��Ks�P��ޙ���a.�`���Y�<��U{-J���*ނ��}F(��r4� I���-��\W�V�0OE6j������/��l�oO��q4���m}���J��ʞ8����:���,q<R�ZI��P߈B���4�4o��>���PX�4Ԥ WL���J;"��~�:�9���
�٢�#��Op���Y@���<)�z��y<�ٵǪЯt|܎��Q`�+�^�c"8JP���*yBӮ ���vi;Hp��&Zu��$�2h�4e�u��&1Z'S�wH���x�_�:�?��s��LH��|Dv2�N��ʼ�B�p;s�e�,�C:���ɒ�ᄁK���R�+!���>���H�.���gr,������o�֠���
��SMy`����^�j�[�� ^�=�D9�DN�믑�Hexk����a��Mf��0���)�$r�_�|�N����_ Y\u_FT	/�[�⛌��c)\��,˼٧�)ұs��|��>C��T��������9<ҋ|��GKx��(���-�Q�q<�@��%��(�7�ց�KS�t�jɬ�k����Qc���4D+�_�z옞X��H��0%G�!�ܠѽ(��+5�F(A�'4�aG��b�!	r��\�"h��2La���݅�+�'M蚈��3\l�O�h�mdS}i��9B��Ʋ_�0��)�hN5��eƄ�pN8�;�@v�gMo��x��~1e�27c(����<�w�2MS�? �;��:�cjn�Q�j��e�#��젧3Bj��YU�����6�[b�/��#g��T�/��̕�s<r�{.��pn����zε�<R
/g���F�)E����D9씇	\3Z
iæ�1���P�ۆ(j�*:���{�&��=�h�C*�\c\�G��:�<�`�46By*{镡��x�����b2����0"�V~R{B��Y��%�0�He�@%,Ďo �#�͞�@��efrS3Ќ*4&ܦ����Zv}Oh�4�|H�t2 }5w|���f�p������+������q����燫c���]�}�(�o��Ʋ�����~9�^��r��{ޔ�;���(�ꨓe�XM�17��AU�F-��K���|�ɛ{(�O�o�Q\	We�˃{x�&� ��t���1�:`�1�o.�mQ�g�Ƹ'X��F�]w�F�)��z59�@�����?i�!d[7�?\z�|OZ �,Z*�*���_`}�GQ�gt���L��H�OT-ʫ����<�x��a�� �lA��q�\D�Æ���8k��gLQ�5��������Xf��&�u ��x��C��I⎲r�xW.=߳6��B�wZ����E�tj�ߔg�M'�S��[���
�GU"n��z��0i��a�;GM��U�d�U�f8�����(˟��j�Q�6���R.��?�b)g ѸJn\Rx��s�څ-��r��ʦL+W�iA3_�����vDˑ2�I��^�Djȷ|�A�D��p^��2k���[7�s�9'g\����k[,Ux�qV�k�]���p7x�'��Wx �1ͧ���P��g�VB�Y��,X}�ћT}.��1���@�x�<[���9x��3p�&2��
���/��9�����.���i��_�h��L%by8�b'b��3�w�mi�@7�:a�":����g�T����B o4��������Ӣ}��yG�l����T�L2��/�ӻ�Jt2���FZ�Sd��iC<4��A�C��'�
Z�]U�7��h�����,S�����}qQ���H�]W,��y6�R�mɪ�Ko�[�f8u��2(z���]��n�e]b��Y�!gza�G�J	�B�o�8����-.�}2S��)X���6�X��w�f q����vx�TV�a����E�A�QWk�DV �v.>&CFsk��t���/�!�ǋ�d��<$4b��c�=>)�M�+�|��B����w�xl��ɮ�J���p]hÕ�q.�� m[�����/z<o�{�X����Pu�q� ��վ.KS�<�/�Q1��P�k�4��n�G���!M���&q��u(QSO�A�n�o��5�뚡�vf&L3�z�81���vڧ>�f::�>����VPݸ���l;n[�8����JI��w�2��
0��Y������X{C��62��:���@�d��2��؂�$�L��Xa��V�Z%��h��X��l�h/���8��*��YP2~.���F_*KQ#�v�{U��,6�q��x��#Nj6Wy�K7q��xP��|�7���1nD����b��;���'�;M�Z����Y�u#���_ڴV�7�bk�Ê�`������ݪ�R�٭�C|�+q]k�5Dv	]iD�(��)��� �2K�(�(�c~ǀd�V���ȹ4ۗX8 �!�㒄���uz g�^U�9�r�f2�mC$!=[��A����RG� $M�����k�.g����j$����&J!�����Pt1G/�߳yͲ��<7����`�Ĭ�.e�M�������zzV��	�����9������w�|��޷+��L���+.��UBW�Zbհ�Bfe�@.�:Ї���<f�:Ԅ|���=kԾ�^�rjq;j�ӊӅU���OVU��=�y��~��S�VT�������!���lƾ��^��e�I3+�����j,@Br�Hx�Y�B���<��pu6Z7%\E��K��G���J�\l[!��Y�q�4s�3�閩���]zdy��"��t��K\	�/�ٰu�6}&L�T��������Vxu��"ʒ�ȧ�M[[���l�tl���7φ",�u�T�8S�#<�NQ2����h��aﵓ�.U����v?.�܇�|���{:��ƪ�����9��1�"}��Ǉ�j[)��}�P�l[E�m�� _�(g����{��p�г#������$«C�X��PT��3��.���\�cT-
�2���T�:A�83"!������ۥd��(^jCqP�Q%k�� 6������t+�^�q��%�?�.��/k&�w���*F��h	����a-��s�t�K�@k>r'V���&����LΖ|<X��1�:���^���t�����:=+t�)>��)�?r%l�7�"�[ʤ�;0	��Oe�I�b�δ�)���#��V���lp@2�	�x�г[���5��&�n�~�|�)��pa|�6Ͻhg�X{�(�x���T�-}"F$�#~�0�������� ���g�e�|'H���MT��'����v����@x�v��������f��ō��ߘ;,�t�
�Q�àysr������jb�b�� ��f%�\�R����ˌ��|F/_`8��(�࿛[s��01�y����<���"6�Y���!��1}���,�� �V�f?4����(ҹ�t�<H�j5�`dɣ����2�Y2���7#e�<���K�&��#�F���za-L��82$c<E�h�7�9�Bx���?�U'�u�]�5P��d,G2�cdB��y5U�~����*0&x9���� ���1��P�q��T��;��K���Q�[>�IF��	����V�ܪ�@�~�{�!o�� ��@t�w` �U@	�:�p�^-�oTYU�*�w�	����J�v��2�	:{���n�3�O�����U�bJn�V���'G��>p�*>�g�����ljof,&�=�1֋��ɴG=�6]5ΫB���b������;f�����Hs)&�?֢b���}h�l�����w�����l���8�@l�^���]̒�F;7w</�噗>�@�X�Ll�lf�ś�E�������%�a��g���&>l�ZWm���$����3�A`q�o�ݑ�W�?�9�\���T�v�
,je�C���/7�G�Q[�
k��4�J�i��D&л�1w{ʏpH���oʛ�����C��y�
X�mW�a�O���\��A�d�k���1�˜��
����{ڈ4����.��'��J+Noh��<��+���;���(d��L�v�̷��� ���� +�}�/����2�����d�Y�
Sf6�j�{}S�j��]K����G���+k8�z�UKGθ�b�Kޡϩ�'^�v3�\L$��e!�p�.�H�6-�-��Y�jX:�t��_M���^��S��;F`����N��V����J�S�M<ڥ���Hޝ/-�OQżn	Bw��hp�`4��K�&��K�m�=l�$2�U������ �ve��m_#�F�N�Y0��b�~��%�5�)<Wr�������Bb�V�5W�)'�[�z�����뾉lO,MG���|4T�Q N�2���9FY4)��Q���?�N;��#�L��N�O��F�m_���|x����Wg7�5��.�)�+E�0·���[��vղ�Dvg�鲮�f��/�2|��`������kû�6cua��DM6^�h��Ć�i4��Q1 SVϨ|4�y�~��8����c���|C���3:֏P�}�0q@Ѱ��Co����n-�`��h�ծ���~��I7��2��� �}oӶl��3ys�f�O������8~o�Е��G��{�ͦC"W�h���$.M?�ɔ+��q���A��x�|�8ɷ�y�7�/�O�� ��I�~��lcx�K�������Z�?7��c�<���F�q�n����|�Hg�>�N�/���g����>U�H¡�c��#|�GN���*ۏ�sV�rc	��������@.dE>�C>@��8�(9����e3vi�s'Ik"^�|z��v�땒J��Z#��مKYG��,�=מ����f�ih��V�M1!��
����I��m����
�s����'�NzU���׸���r�6�3�=Y��0�4�܇՝�l��nR~�Oo+�4 �Ѷ�Ѯ�fHiT����S�pg��` �hL1>dȹ*A�:�crE{�Ǫ��\/��d�zIym�4C�9V.�|]=T��~ �45�0��gJ���®p�����/3G�D;<Q ;	�3c�>���j�b��&���Q\�- ��� R������_�ю�E���G��欉<�]-��)�Q[�j�L�>Rcqʈ4�1
��9��p;u�<��g���Ο�08H�F�t�^m�Z�Q�K:�u����VPБ�HX�#!f�hZ!F�'z�3p{��a*������P�_����;�{:D��Y�t��Ȧ��Ӭ�7VP�F�{q5�)�yUt~���-��r8�\�S���	�'K$�C0�7��E��Dh���ۭO8%T���jԛ�v1*��?���G��X�^H�K^��ǠLJ�GVX��bk[��:�8���Uj�v2�E��A��&L�;���1�Ҧ��/�`+aE��@�"r�B$i�����7P:t�_�{C��u�R9���	�Q���� �s�̫ɲOٕ��F|�/L{������G�I�}6 _/1Q���@I^�v?)�o�2�M>0`j�A��T��k�;��2�?�W =����Թbz
������V�c&q ���d̸�}]�a�B�{!�qp\��af�č&��>�p���w��x>�������H�r_s�p��l$��`���H�MN�ݜ�I4$�ڔ�M	��8�K[%�����j�w��ֶ!*Z�ʃ��� �=�������@
 ��FZr�:y��/{`%a��Q��,;95���Y���zc6����R'��5�2Iwp啴�M�r����3@���ȸ�ͮ�0�H�%�42�ά&�����'�1N�Ud�0�Z���_{N⓵�]�9��hhe�צ�O��ѐ|��d�J�(g>3�)��q��'T϶��_ln��{����վd.^��O_��W~���hߢͫ���XBiC�3ai�Uo�C��n�x\^���Z�ӕ �4,<5oi�����2�#h-b�Y3>C��pG&����c0�Z�_���H�H������9zt�vj�����4Vu�!�)����إ�62����K旋J��[������w�Y�v���WO��3$�P7!m
���q��A�n�� �:��I����kx˴Ԭ�o���:�C\�L�7�������
�X�E����������_A>qu�9	�dǑ�L�[$��Ѣ���3�c\�-�[ ��#��GfU+ۉ����`]��(�)�A��F���5|X���$�m>*�t%�M��-�*��X,i ^(���˶����_����ԙ"��y����iM�/�B���xJk�h�Ƕ�i�u˲6{����8�my;�j�{JK��L8�)?����Nt�Iwx�W��zy8���WMd$˝7;���J1�x�b����Ss�k���z�4�50b�h����`��{��l�nt�l�T�O�����׆P����3o��̳�&:ϥ�7-X������(�0�7�\�n���oˏ?޵pX��2̓��1������k�Fs�BK���������g��}�l��b���'�'B�p�.�,I_%�JK^{�M^DK)*m�F��d��H�k����Je��vÑi�<��#g,�đ�4��K�AkF.���\���ps�suA|�< F������$V����p�+�G�j������ �B��s�ӳ��s�Y��p�l{�z|�r��}�M�3_�_����:c9�mߋG�͏�0~ݧ����Q��`���K(�/_���s�V��)��+��mmH���k"{���=�3i	a>e��)D��Q�M�ޒ�����;������&랝���q'ar�MCE� C���TK�8A�	�$<U��֥��xB�#޸,~C���
D��M��qgϧ@/����*v�� 
����F�%-�R�����M+F��矙��[��NK=��o1:ت1����^.�����Nvg�C*�riI��<¨�P��W\.�--���h����}���9��ˡb��-�'L!a�F\�x(�$�0,\vF� �5�xDd��Ej���t/�o^FuFR0���U*���Iò��;���Blf^Ɛ�A����	]򒮤4�2%[F=(��!��h��V�g��=_w���S��Q��/�K8Z,���{t1�h���;4<����"�('K���G+�BS~z�y�,RP��`lěz!P�O��P��m\��y�0�<+g{�����C��)JR���.E���k?/Co�N����	��rN�;.����� #-���WV�y
��#<aE6�O$���(㞂�ÆJ[j�6�,}�`.�PprD��0g���R��!;��q��#��W[e���{�%V'�h��j4[�՜%�����W����X�%	�w��T�5�-���O�&ggw52y����Z|G��8��l���<�#9�Keo}�﨧�*[�� 1u�ocbE��vұpиO��R�]	k{~k�!����۟ShA*�\�;_VI��!�pg�YM�5��B�fc � (c�9����˥��R��]lx��ᖉ/]-�`������>�qy�ҍ� L����zsb����yub�����UMX˂��q;�)�>�-��',Ld<l+/L��B�-n;��56��{O�-a��of@ц�5��g�Y#\aa!�6U$z�N�hBecB�$x5xȊ�iO�f)AD��Z�Z��Q�h���.v�	����g�\���;Z�@���d�͟�CJd0܉5�ZߐK�~��V��K:��ٸ���As�}�ף�h����B��ъ�E��ȼ��"�#�����;O��� ��Kx�ʭK ��p�D�	�m����F��|�LF|JW����?��	t��{L�JEp�+i��F�������7���@��b^ �C*6!���\�����7c�!��n�������.�t��bIO/�c6�f���B�������	�䎞��kQSF���ݸ�2=?I�]2��;���ȟ�H6�_����� 0�ѓ:����/J������2��J���HރCiN3~O187��.+��?|�xi^�_o�\R�x���&��)-vY��� �nwy��Vз ��<p��g����N	�O^IE�[�d%�^#C��[�&B���iu����ų��V�7����n"��2t�T[j���ĵ�X�w#�u���WU�Ov�]���Im�
�1p�c� ���`ҍ]�ʚ�*�e#s�r�v��.췡9)4��-��#��ƥuֳ�>��1Y�&m``T|T1�V;����sg�z;��9E���V>�+J��m˖�c;N=%�a���&)\����neqvX;{O.�������u�>=��qF��5���0b
����B��~�ب�k����R֏-m����X1��?��/BΤ��jj����6^:��MmG�C�,��֊�H���j�n������>��<�8;�����B��:��qn����
R%oG;OQ	�{�Bc�IjMZ1���ЯGHV�h.�YX�=��)q�t�L#�m}�K;]����Q�2��-�������n5���C�{C���S�!Yd�Cv0�{Mi��4,����߁`�2a�XJ礑�Z���QPM}��0xJ���P�p�ϕn��$�ub|x�=t��T:<�[B/�h��#���pV��s>E߆�"�B������o��EN�]�j��~���\��������M�[��P3�Ve2^�:V�Ψ?U6��	�������3@bi��%_��X�h� ��M���M�9�A�6d�9�������>�2ф4��,��\�y�T����$΀���8�L��b���N�D���Kzp׌\K����b�Âà\��!��L��bfYc���ImBL�������a\��D��@�f� "�FՃ�8Fx l[���o���b�kh�)(G�f_�ĝM;ߥQ|�Ez��4G��>�5�U%Em�?D��|4�. o&�cF���?��4��W;ߗ�O��u|l��5���[���H���+�MV�w�W�]M���\�v�?��zX[���V%��+�
�nWf$,�� �+�skE��of�-�{��.o�H"����og0�w���~��`����o?�j�SĢ�=\4|�b��R�H��� ��ZCC&8�M�/v"L�N��p��j�������;�n(Z���Z�4^��,�D�������!�:aʛ��.�m�g^�3䤀@��.Rt�4A�<�_=�a�bQb�����՞�$+����X������
Z0�:J^�?��ጃp`�?7�B�ʮ�@*��> i���$H��>��/�)~1�3�1ee]/���z�<���k۹ܔ�v���^߆gh����}��o$M�ˬJ	�j��������*��,YZ
,QW4縤b�0Wɡ$	c�;N�,�oe8F�bR�@���T���¦�_�l>	Y.��r�)L���"�U����J�h�+uh~���t�sG-��[	��!���ek1���)ID��Ț;<#��M�8�PS�2�lR?�%��`lpMq4�<��Q���#�O�h�RI�L��0Q}ʰ$y�j���F'�/�ۅR�p�&��jk�+�"_OUQ*ل�esKqph	/�l����C��%��q��#��pD��贬��K!m�?p�v��,�C(����������,�����Ｄ�ã[��喟��r0(��ZK��X�U�pd��s�w��ČV$8�\.V�wkOv��s�i<�Û��+�9�/�x�D� �g��:U]6Ⴢ,�= ���Of�~Mݼ��U0��[��CKD.N���{�ys���@�� �X�l�-�Q����'D���VL픒\���B�R�������y�/z�͢A��m�yY~�:@{��N���),E�Z�����RO�P�rQ�l�����d	�2�iD(��LW�֞��%:IN����}>D�6����9��/K͸v�*#(��Q��Nu��Z���˕Ѵ��g2-��ik�|��K~=�<��/u�^�� =�a?��&�T��,�jc�8,b��S�|7.�o3I�G��3L�ܚ�w
!�\>D�e���'H�����> �Čz�SS���k�8��RA_�h��0�J�����K$pz�G��\�)���w9 ��sY�w�˘)�0�#����0���5�rkS��6>��#�4�߲���ݴ0"��w��x�����!!���f���6���xx�.}�Ħ�ZE)�����Mk�:��j���b��Yp���-eKw��Iq{ߤ?���A��uṿ-��%q�vWC��J�h�_q�As�Z$�߾�2㖅�v
�1`�t3�ي��XZOG���z�9�q�ӱ� ���$m1�d8����kǝUq8���S�ÕR�D۫��-%��RR���� �L�;+�����_�Ҍ=^�9Uֹ�*| ��ΐ�=���:�R�6N�^e�1�>��Q�G&�T��%�O�U��q�"�C��۹Z^���Z��Z�"���E@_�V	���Dy��]��뽤"��?ƿ6E��*2��Vz�n�����9���g�g�(=̌�^��3WH[	��_�K難�#���Ms�R�^���z������}U!�U_*ƴ6�ʦ;����<d1��,x�E�要�795i�w[5`@!m~���v��f%*�}���Q�����um:�ԢB>�u��y~gzA���?N4�hF�Ү<F����]��#f�T�`���u�$�/Dwab��E�#�k�����
�1܏������-(i�UÄ���,���  <:2�P����9k��g\�����d�-4F�7�1�W����y�w����P憊qPw����n���ek`�n΂=���0W9�A���T7�.�q�S%?T�q�j�/e�o�ԴS��ۑށ��Q�O�+4ȁ�3q�_Yk.F �ױR�{��h�ye<�Q�@8����3�u����$��M2�?o6�=1۾.]`�����,<�ӊI���?����b��䓅'��A>5��[�D�N�� 0b����+�����Ax.o���x�UO1��|Ɣ`� IO�_���h�U]�r����9�-3�(0�t(4� n� �[IA�4��bՠ0 sD���g��I*C_@L��G��h,�uf�nr]�|�O:�o&Vvr3��̑ш+�,����Z��ť���
��N'/�Ijb�+Wv#���e-~X�n�8��m�[�Nxtk��zq��'�s��Jw*7��D���j��!d����Q�4��BQ�1�<.+��HѠ}Izdm��Q��%�nV�W���=�<Re�0'U޵y��6�A��.��^r.";��"����G�SwM��tP4XX�BQ�'3X����!��[�Lb���^��w��6�3�� ����J��~���a
3Q���JU8�WzuA�uv�ջ��Uxc~��}�O� �Y*;8�9b3�3�ڬ���aT��<M�
���=G{V���U���~<s�5*+Iº���w"���N�UhA<�u��e��w����٢��[�U���v�˰�@>l2"Y��J ����Sm����^�3���.�/#�*�x��
�?-�4ϦUq�ι�ث����eC����T�B�m��H�����B���_������2���Na��ώïnD��S����vNo��(��d�����5�^�tUQf'�ƌ{��l�Ue;�	O`�I�����K:ÖJf��6�p[��M0�i_m{���W�䅪w��Wa6�P�%����h&)I��
������ӚSe90���
�`�����{�p���w`��9"h�K��~�8��ȭz�5���"�Z�KV���$�7P&���{~���ʋ9`�Q'��8T���X���|bb�mi�7�0�
	�.���6�A�L2���� 3�eœ���L<niFH�.	;6���w���g'�#>�z�Ҷ�������L\*��FF*k�/�����^��U(��G������W�}�q�p�REj�ܶ쉞j&wK.��ocZ���0�Bq�2~X)E��1�Õ���Y�[�QSO�o���Ck�2Wf�1L�����<�z�F��6B�l{(h���K9,��u/�+���<R��b\�G�aV@̧�T���p�8E(
�2~�r�Yqp�U���U\�$�$�JifÙ;�I�s��YHtVK(��KǸ��)]�B ���R{=Z!W�*� ���5�j�j�p��S
\��� Ⴏ;�;�m$*gb�A��̆�����Q7�v�JĀ{`/"e�r�ܕ:k��KE��;Q�yv�*�y��4�;��^N�Ec��`��%>&:�4�i���4����w:�����;aKN�0~>�	�w��D�QwBf'� *1�����<�Y>HB)����jK�Ԍ}*m�&���!;h�̒`_����Q9��f'iBeIz\ˉ�y�z������܉u$�B��h�07���Of�IE�'�ˣP���b��Hw�ܝ�!���k�ҕP]��A�֬�D�����1d8��lT;�J�qf@�>\xBmQ���@X�$R��]0"��K�q2�I���x=kFt��u�&�ea��Y-��@�7Q*A ��8����Q�W��_b��p�-d*�;I����!6�k<����-nzN�/n~;=Qp�<�U/[W�b�ſA(Բ"	�8��3o,A�dJ��fo�q��0{��s����'ҍ���W�D���j�K��L�q;�u�܃Dxo�q�=�^QgT�"@> �g��xI�b�,�����J�*kU틂R�\���ы�ɌP��ӟKκS�-ˠ+F��I�<��&s�Q���s��l�y�~��83�A]JT� �e���[Qm���}���t<����>��]��L6�(��hqK ��rӯϘ�GK߰˝O�&?��:爀=[���?8 ��3{��Η������x��ˀ�Nq��+*D>�zLY�Vu?��d:�T�~J���9XDwdV$gE�;#!3g����Tum�9���H��q�iYIu�%*D�㵅`ݥ�r�BF����3w\:s*;t��
��.����3c�J��G2?-�9���z�E-3�u���`P�G��ܧ����e����}�ϙPT�A���-��m��	���l�~N�˖q�dN�ҽ�,B �=������c��'���%��>�
t�9�5Q�0n�S����������-%-�ϡ��Hq(|��G��2������y��Iy(�Uz6�y�5s��q�YY/�B���m����}������#U2��Gg)#N��|��ya�+!U�]]�3�NO�r��}՞,\z����!��J�!m�.���.f*u��}f�gz�ŷĻ[kI���G�XZ�ʂ)�])�[�uU�B����v���8��@{^�%ϒo0+���G�|�y�F�+dI(�ܖ��zs⍿���!Px4�0��\37���ۛ'�2)E^K�	l&�C�P-�0[휇�}9y�b>U�خ�#��[E!_��F&��w�E��.DL˿#4�:�����&n�lρB��x���񒃢V���sƊ����"/��~��8I�M�-�JV9��x\`����9�)����J /'�F�W4i�wdd�������b�3k�~r!�Ap��6�{F� �>�^�;񻨓/����uHSOD��!j�$MKm�H����-����S�;b%&�@C���s!��8�!6Ǟ^k��������[�ёcGi���t�JV~3�k�*T��"��X��.-t�L�Hvh8Ϫ��{6�o��V^� ��5�3��^�.��(�}]�����1k#� �K��	F�.e��qoU��r*
l��QP���i ���M���1'x*,'{(�/p`�2K��~i[HZ��)��|a����Ԭ�%��K[Sw_ce�R���:��2����d�ͩ�-��X�+/v�NX�Ӎ���@j�Jr�|*{�֤n1�_4WF���"u�K��y��33ݰ���R�Y�Q���L=1��T����B������	y-�}���&٦q�]	�G�]fC�#6��R�kI�ص�0M#\X=�HQɾ/��0K�/��W ��1�E���6��-�����X۸��ZT�q���
���Җ��^�ui��7W����J����u�W�s�[���s���5ͼ�{�a��8�s� ���!�2���C�R e����H75�|4�b��l�H"_����ڭ|���f�7�	H�u�5�B8��]�sl[6���q�/F�P�x$b�06weҨ��n�)�;���k`������J��	.����оY�ɦOw~�W;¼�U.CI7�����l��t5\3n�oD+l�j�]�p�{0FQ?`�&^����~ t^�5�
��JT�K#�f�rsoF�'�w�
H���}�h�P,	�xg�k��ߠ�}w��]�p&��Z�C��J�Tf=8�rBu���_߈�c���3R�S��H/�RX������n��Ks)��:��!�DZ�O��S��Sv��rce:��I��o���p���o�g��41�A�R(e���F�7���U�u^���d�����S�O��r�
�z�	~
�3w`�:a���E����T�&�<Hv'�4����(_ucChW:;B<�o9�,ٵ���Sנ��;j���d��Qa#fR�5��`�>�
�0���%(�	�r)S<�L�4��?�V\U���~n�mB	��o���6�R������4;	��0� ��5@��#["��>�Z累��5)��|k�N�����H����{�d�U���v���RQT[S@��"��(4x��Lgg�pJ����,E�:[�G������H�	qP�ߐm��EkE�˃�
/S{4a�!V# lJ�o*m&�Q�>�.J�k'}�2J�߄0��7�Ѐ!Z2�YMn��^����w��[ �g.�����u��#��KN��D%�ըi�d��Sc�<��vji\n4(�}Q4Z�=_e'������c�������zQ��t$Мpǲ�>$i#~�*ZP����-�u����~ܗ�5�P�uC�g*͎Gc�� �<��9��E��������c�������G�b�[32�^�\��V	�[%��K)�T]���}"��_�lO-I�����w��܏��y���Ѩ�i{������i��7dժ��/�R��$\���ƻ�8%
��H˻Cɻ��/Z�ٛ<*�ӆ��]��	�c+?�2�j�@�D��5�uIqۃ�bَ�r%�RrˊåP�����&qn�;�����bZ��خt�U���\�1���w��N5兜P�|����P���1vR#�`\a(��,w���b5����ᩁ4��gs��L2�^�V��Fa����w��*���d��p�[TxW���{B� �߿��U51�^�L.�ZR.ޑI���Ys�?�#i������ ���)�;��T���Z��K\S<]m�n'��l����r��G<�,�vB�͍��l��t���_~p�Z�o ג�K���jĞ�5.�!�x���ngmG3*kmqk�t�={�}	�_�3 �3kt�����ko��d`*�.>*C�&��OyVQ�c{��H������9�W|�z��ym5�m3�>�Kg��č�Zr��VW���#X�R_c�	� #8��XT�Ga����8���l�_Oc��I=��={�t#���~GAI|�
}}ña��e#o\]��t��f�z�Ë���`�/��i~��98AO��aVMm��[ic�.vE���)~��˻�[�?YxAG+�En�h	���~��Ч�ڜ;����в�!�q�v�eQܭ�`�N�R>�QbT�E�{��f 1G�n^�yS��ak��������:#�#c6),&mM�y���C��r�M��6��R>1bs�=[�V���6��$N;�� '�Tal�z~�)I�!�̥��W�ɦ��X/K���㰒}���O�}"`�-J�M+�A,���J���x�s��Tx6ⅈT��w�j�q6�|w����dn��i��<���	f�VC�˄<]>,��y'�=���<ڟg�a�l��Ɗ=D$c��s�ɬ��;��!�l�^��d�!<G��|��U2j�pn�;m�!����_ũ bN�g���*�x��BC����7�~ʓci��,���*�s��E*���OU�y�>$za����Ú�Q]{��e�(��Kj6'���Ƚ�Cu\�|qg89v�~R\�R\��W=z]��9�m5��r/�ĺ���!oK;� ;���g$��8K�͈���W
�#Ga&���>+��lYx^_�(�IZ����@����a��vLa��$�0�Y#��D�#(Otן�/(�C��)8SSd�߷�[b!������>���r��RZr���-욲�AGJ=m7��_��`f%�um�1f����@��,hPµ�U���俲�% �;�
Y��V��J�}Zws\�}?�C`̼�����h��2�X>2��~��nIoK 8��)������xfЛ��ؚ��9�UNY�d�����P��nў� �⿆I��������<f�U ��6 �&��,�G.��w��hh6?��!����q���Z�l��Z�ϫyj�?��#1��
(A���|�Tፕhee\i4<`',.��y%�^�?'�Ő�Y��� 
��9>ÿ�����/�q	s��|�u�L��g�s�����x>�x��{h�-/r0��E�iW=ٞH���DNv,A�g��#h��q�$�"�:�����Gu�������v��_���7hh<�~1Q��I��S�D���&<=��r��e*�_�d����}p�$�׽�B0�����9:�X#*%�t��pگV}5�S]���AY��@�X�����+�V�]���[f���2�d8+�=��r�'��S`p�����N�)��v���q��lt��l��'����q�%�)}hZ������k���ҫ�E%�c��!�s��5S�/�D���
�KN5�V'� ���� � ���Zi�6�51S�}�4$Ut���MϓA~�3��c�2�Q�����L�븀D�j$��Y�S]>N�ϟHF�N��/-6h�L��G��hT������4�VEq99��N_-�]�D\~�d�ӹ��d\N]����V��fU�@�Y����1]NY��=��X��TŁ���a^]fyW�\l0��F��L�4}n�(���t�·��0�-�-���^]��jEő�HㄽrJ����M?�����=��_@'�ҋd������Hk���&�'k���=�ܓ
�U�0�܁A���c�[��O�����qK�P�����PN�J���H��PM%�`��Xy��������z��@~�ƫB3jU�q�Lm�[Y�&*c�I���Bҥ�~����U�%�P��4.�q�*#�嶚�}~���(����$��hI�=�C�ar��g��i���bh��c�yG���àA8��>�����ɫh����9yb	:����M��ISv23&ْ���<a�Ӓ��2��"���Q}�׊"��������]��k5�2���?u�i��JQq�	Mw�񕼧�����<���_�$��S�yE&��iD*M��&$y?U��X��A;���Wu��vӮ�l$G���R�v�ҷ��b�t��}�@	4��9cO�67w�Ibe��)�J~ȎC`8!hq�.y�t�Q�P����k����1~
�<��j�F�L5������k�V���\f�'^RG��9���\��v^;���&O����U5�e�6H3�p��L��|���Jr����C�1���n��"�veqH�����{���R�M]Șe]��:�C��W�ȍ횑���]0��d�ɔ���
��"/@�g.��0K�e�1R];�z��I����VNYZ��P�q�v�$B5?�	�ΎPێ�@��9 e��À
r�9�����2@��\}w���-��[*�l�S�7�h1B���ҽrhQ}1�Zo'�g�?	�I�{p������X8���M�VD�͑��R��:��V0�CN�ef*���a�ó{��_FoҲl�J�.�.���_�v�Ӓ�W*�g�h���r+z��:e��J��1�)!�/M�����d�ݯ�v�m��f�OO����2vʦ)')fT�eG]�,x��.h�Z����B�c��и|9b
�Ss�E���ѻ�?��c+:��2�ؕ�L�򅦭t�6�a�a������d��?pW�d�A%˯�ɮ�qf�����%5�'�_2�O�V����.,k>�� �dг۝ . +��Ʈn��ạx����6���k��AW��&�B�����G���Ưp}*�<�T�D�>�[����A�c_���B�cy���}�b�!��Ѿ:�+�j<�nlO`���ϸ��Q�*�����epT�IA�� ��{���c��:l9(T>������41<;�_P��U� �*h��1C܃���@�y'j�Y�T�YF���`���6U�l���2���m���M��HSݲ����VÁK��t�v(��PwW���¡�[v��#'�d]m�a��Wv�g�&{�te$���hi-Ò1�})ԉ0�x�'ƈ�>��i��S黛���I+"j�1��-)LG��sr��t��0��a�A�`&��� �G!tBZѲ��o�@ت��<���D�'�#3��ш��I�=�M�MM���ҋ}}|��{X�O/jJ�=Lw��~a���WJ�����2�<C"~tn�P`n���O��Ȑ��B^�p�ǉ�ՙ�Ed`B�C��0"�@,��eT�ow����apB��B��Ni����i��j��
f���S�|u�J�7͡Ƨ�@�2�����I$�{V�3Q��׫l�6Φ+�|��s�����k�����/��o�һ���1ȸ	��M��BJWL'�f���T(�רLer�b0��a���C[����p:��1�n�9U���Z�,7Q��kNzRZr�Ђ[��nS8����'IQ�BÇ��qj�F�}ȃ��{Hp��IH/M�:��`g�R�h��MI��&�(�7�Q'�px��ൔԆ��9�ɨ0�)�#W.�v��Vl�ʝQ?��
�?�$�xƔ�*���`c��9�G4Et������9�=���إ��.����Dr��X"�_U.m'�9Ґ;����������Sov�G��ĆѺ���e�{������ֵ�6�K!�� ���j�W��g�XD�0��(�O�PS�lTW��� �in�h _e]�q���J
��Z�
�#���o��~��[(_����RV����s����FA���b�9:iGe������L�IOL�_�#�_�,VQ�EW���l��A�v���Nw
�1�hp3�q��/�� �� ��=ˆ����(����� ��l�I9� �j�;t���9�CS�<X��-FA=�	�9)cRT����~�i��w>m�c��U��F,.�>X^^���\��Ŝ¥�T�sb`X&��3�^$��#BaհP��,m�#XT����o��ǘ���e	~r�sH$��&�R}��'\�Nf�\�cO��T(�K ��L��hޢXՀ�F��j 9�w�j��~���	�0Y�	T�A2 �0��}������-�)�O�qK�]��f��V���*��v(�+�rcP����	��y��_8�*�Ә����+x�I�ĵ��"��&]!��������܃2�b��쩵��O��{�z�k����?�!H�{\�w�T��!�]G��j���9Qi�"q� _R�0|Ǌ�Ց��^�}g~v���%��U��%.�V�%���Ic�W��W��ӷ�� ���Q�m��e"���u2���
�6*>ү�(�N��Whj-,X	�\0'D�e�L>�<�f����B�gD�&�r3���v�쾇8��B���A=F7$N�~,�@:4;�e�wt+~�E�*�	��-W�D1�9��t$W�W��	��Bl5vr���Γ���$)�8*��fA������w��>XQVi�F��m�`��e$���� 4WC��Ľ���Ư�
.S�\z�8�;B�&"�Z�J�^Z~��|6�ف/#���/a�b��p~r���i��-\�S)3���q)��\W�x]c��c4���̪U��/��%�w���}>�c�f˼��W�e9?!�G0!F���Q��&h�߃�S~X����и����<��G�2��K��)��gڥ�B
(�Gx�r�x�6 L��6[����s3�����k�ְ�!]ƨ�.�X��0ƬH"���.�퍱�N!)�k��/�� ��C颀^ ��о>t�H+eފ����l�́��)�S��y�6��׌�/~�xք�9����d�Iyz�'�"�jb�o1f�]܌yQ~y�����l��Qn�O�WD�㪷B弁n+ބ/�m��2�J��)�2�#��~�Ue�e��7pU�"������f���A q��H�y�_q2g��|��H��T�l(}����Z��v�}����}�:?�_~����,S�m�.�[tіX���� � >gw ��ԝr�����e4ێ ��T}��MC?�����'�@I�m�[u��Ҝ���9]��Xs�%9�N���v��<S�<}���"�r�	���ڈ5�W�S}�_ihN�;���Zn�a���W����"�j��F2]�:��%��l���ܣ�/d2��n�w8��ek)�/����x�<��'���l�J�s@���S�E�jؽ%m1�$�s�<D��T�j$���>�+]�k�[��D�4�J���E�4M�uf�fo��z>���
g�7����ۻ�dLN�ɠQ�[o������B���,\󅬝ˠɬ��	3��+���\�x��i)y��[0��^G��>!�:zn�
��*����6J)a� }
���M@l�
��u�ߋ��y�|Rjn]�1�јQ�������Y"�>Q.=�`�ǉ�?�X�ϔ��4hDwN��1fXsp1u���1�.<��<�O�cM\p7�EIo2I��1�SJ�����S��#f� �2ح#D*>�����1�T�|���Z����Dʩ�@�K�E�"]���ݶ��~H�Z��R�l��E
��w U����h��^��=�Ƀڿѧ�w�C��|n�����1l�.ɲ9NeTPl^th5F�EraJZ ��W)*{��}4S�}���v�9!��F�J��T������>S�q�.uL�|����U�v�������o|�7G�)�
��h�� Ȫ�����V�]@����Eq@�\��DR�*�֛�4P���;$l����$����o@�m�~��p�^���!�%N�������<�P2��ֽ5.��>a���$���z`(]�Bb���}�ZE�*6j�@y���7�M�����N�gT{��(��4nX�[ }(��4=t��q8�H�A����J��5Y����{`���u4fZ��n��_��6��4U��}A�i�^��W(���+c{<�\�=1��5���=�rR\�*-��p�ϔ�����i'YgW������dܩ��9��*�cT���G��%���c*?aU�z���n��7�3�bG��c���*8Z��T1�E���F�n����R�!��2b?�!	�+�\m�f���w�~�;a-0��ol$b�w�BԔ� �_�����Z%֠𙻢1�}n��Lz����3�C�2��Q��ae�����>�H�?8)�;�=~WSBw�Ɛ�S����#�ސͅ`�i�؋�p�(v.�m4��iE��+8�Z�����y���_��eR�ȷ���R�������
�%F]h�+��@hDp~�t�\9;�\�+������)�xJ8Roa�R�� �`>����t.��]���&��7fV!��O�������� ��M5��!C�(�)Z��z��KE �p����iAU�4���'�H띑�0��fҙ��I���~��G�1�����\@�k�^���Cl�}�/�>��?3Fc?�e^��2�|"�(���ihJ��!Gc�v37u�X��S8X�RR�G�=0���!25Z@_.8��&J#��'d�aE˚j��zw��I�E�>�W��[�-��Ӏ���Q��S��5��r�Ŏ��B��jRb��P8� ��3S��F�/�4+��:�&�B��Ln�޺�|�M�S�f�Y�O�|�@x��-._�#r���Dw�n�%��m�:�6���R�f"Jﲌ���ܣ�e�Us�c��0�@9p3>��[�UH�[%h|���j/���$h4�r�4�Gi7�=4R���~z�e.���ה?�}�P��3ҦqӀ��rK�<C�HUh�F�k���:Q{�N*�ޜ�?�F��c���Ӡ�r�c�T�� ddI��}(������� O�9zӀO��>����!c2�nt'4Cl�~3��d�K�u�H�[dn�ZUJ�)�lW8���w���Ig�������R��w��%�����
���zP�I}?�!O,*�v�� �=�mM�9�k�"e8x���ϫ���b:1��l��PwK�F���_�&D�l�Ps��ET&�E�b(��N_�;w)�j(8�$�"��'��8�uϏbJ�Y�\�����p*[����8�'��Y��V���[O��sRsP�s��aL$��߭�@O����~�Q%OZ�3*}������v9x�ݝ����O܏e<�wKJ u�&9.:L����b��D��"�݅X�[��Mmy���\ɍ��vR��G�y����̄�r��,p�p^+C,�)��x��:/P��������F�i���Jj�NA ��X�x
���
��fvW�]�<{ �� ��a ���G�+gk;�u-�9E|򳄰C� �p(X���	���x�Zp��̾~l$��0��dߣ+�s&^bgc���<tQVw��Y,����=���Nn����=6�$v�T�y����A��ٳ�C�7��l����,���c���������ׂ{�,�r�:k�h����f_r�����0a�7�F5$�b���l.	vn�O<�:08R�ܼ���u�BY��֦��`��6�D��5ɾP݉L��l�k�T�[4��/��6%ж��:H�2��2e�٫ ��gI �we�Y$�r1�B�V��'��Yp��R��Oa��Aʛ�'a�t�ݎ���@͌�� ]Gs96Ѧ���iH�rWt6v��!�M'#9��{oT"��ƍ�Jz��,,8i��ԟ}�K��$�o�G���1�����Q���y��ӑsa��}#�����u(�kn7��T5��qm�������Л֑�C�_SݰZa^�L�?6R1�� aMto��Oe�&�I��=�K�&Q񙿠��NQ���4�GՆueb�-yִ1��d���C+ ���C�@��%d'�ya:"Ia����g�M"�b�C3��Q�Z�!~j�C�����y-��؀�;�.���!�xs7b�H-j���Q�C��ҵq����()� -�co��9�]`�A�l˅Z�6�k3�bz���t<}�[`�=x�ȁc����b�OՑƮ_[�F	ɲ3�3{T����;�+�6�ŀ�������+��Alx(�� q�Rfͯѭ���7*��%,�K��d�R�k�>ZL�{R�����I�;a]@�+�­tU?�I����y񾮐�H���X��5�����	_��U�#���֮�vb-��Ղw"�Ua���#e�҂,4�⍂T�SljR�|�f�R?��Gْ2�{`|Vt���``���J�g�p��i�#�� ��n�����}2x���{dxU4V9���4�X�z6�^�frhXГ(矲Ϗ����w?��Jh:wdX��	� ڕ���l�od|ֻ]n��Tͪ���J~J�/�ϡ��4C1���gAʪI�eb��9�f�����hQ�>��1�; �;���wu����gr�$`��?+��֐�x@3F�S��|�.��oUf��h�._xQ��Fݔ!����G@g���s:��N������+y7�]ױ;�Kߞ�RWr̸r�WZz�������*R�g��H�׻�n>X9�!i����6�y�ٕP��WJ�W���BF�CK���%���YF�Xmر��ݨ����P��!<	�W`�:���xU���yNQQ�&Կ|��- ȯ�^6ˣ��W*�~�L��UC�B�1Q�����p"u�V{�&)��F5
"}Z������U��F�H$���k�^N�'N-_�%���Y�Սp���C�
:�2�����M]8k#0\� �cXG��KN�*DX��۽��oz�I�����'~Y��edG��s_:|�x�9���OA�g�;�6��A׀"i����g&ZF�>�W����Yo��;�7>��^��)g�E�&nN���#��Y�%�y+���jN����c�e��H�*�O^�MQ�A���g�~��n�|��CO��+�CA����Q��;��6u���ܻ�r8��?NH�g_c����M�N2�P��̦k�Z��'�N(�PCغ�W5ߖ�L���A��+�3!�b�Mb�L��v��A|�o���UF�S�9/�g ���)��Z����BYI�A��=}�S!r�X�Pz�u�\k���l���������c&�f��h�����k�]�F�)�p�g�[aY^����".�h쑑:� ����Cˠ���1�r�eP%N��Z���c)4sff%��@#0x{������g��ߡ�ndq���LT�1���o2�E��Jł���f��4[���_�C����Fya_� �a�	6��#}p@,UuG��ħj��գ�AI������&�X���� �����Q���u	TE��Q�C+� �?~3��ۃ�Y���M��z	�;
�fI��]8P��p⥀�g[*��p�C(������>��9M���ک`3�L�.1�y�
z��D�s��h��P^k�U�˩<ļ&(��-�b%ñ��$.��pl�w��d`-��橚@�W	)�)����>0�|�pu
�(�N���9;���$����,�+g�u�^�D����A��a���
��0o��<AzTs�YwM֠�0.H���9��z�]a����X㭬�k����2�[;<����FLȿ;�z�F.v޶D~����G-���jd�;�����d��Y��h����n�>'�s����6Y�2Cs!��E���"d��iF�e9���n�kK\�z��V7��S;�ۀDO{���|�Q�$$�&�ll��Y��һ�K��XPW�ƔP���^�`���G���I8�S���,MM�4����ݏ�.���SY`��5��c�n2Y���bA�;jw�X)�����R����uy��zA2��Ο|�������q`Ե���"PwΈ.H
N:V�����
Io'�Dm
��)�ynA2��g'Qh�����Z�-�,p�_��.7��f�M'�g@|.l��Ԝ���O�?wA:�~�],L�k��!�CCX���mޟLڣ���IE�z&���v�ne�B�zѰ�Ş� �|�]�i��,���ve��+M�W`a�A�]�8�gf�$��PO�8w���@�k�c���3��n��\�*^��̽�5.��e�V8�����3������_L4��q�L��Eæ����t[�k��(E��X���;a����DŔ��K&`Ĩ��yx
)	�^�m&��4��W�N�KB�֞�[zAo͇XI�3��㵮,SZ��l�,��~�{J ��C��z�a�ai#Vi���ڢ�[�+8*,@�yTM�Vf��H?Y4�5��Q]0�L��ˬ������X�.�rJ[{�7�\CK	y׍��b�ڼ��S׺\N����.�j]��×A�?�K|8m�&K�,���h����,�x)%�J��!���!�"�v��}�n
�v��j�r�9u�w�0|�Et�u��B	A��{G6T�"�?��0�g�[Y�U�{��w6EH*�P��[����v����W����s���慯\x	���.�x� �#7���$B{���7�_��	�+F�^d�tp�'���[��cd����$ਸ_,#�!��]�-5��&wV׆�'A�2�d.��l7C�ch�r� ��c�ʇ�LΧ�ap���h�6/�Q?�#5��/��/X%����v�w�'HwO�nV��vM[�8@��n����XN�����5��b!7�m�d����#�R\�[ë��c ��Х�����03��\\"�A��m1��wgR��D�a��?s��#?��L��I~b�nݡ�Y$�( �l%)�V�C�&�le�DԠ�r��,ɪ#�/ě�7��/�J�/>wڴ�q�,�(�E9b���'h�k�h��
����S��k3�L d"4�b��xs��w6l�9bҲ"b�NF��X�Sc��X	��L����x��>T4�'�E3])	�bk�%t�J"z1���U����y�p/_�2����/!�N����ؕ��S�N^����l]��2���F�_$"��Q5���y����W�=�Lj���K��M��x�Z��r#��)�>��{�%!y)�@U1X�%S�'�o��x(�{��M�(��F�o�!�R�
�>�0YL(������ؐ?8n�+�$�\C`�';���P�,�:��9�cFڒ'��v CG����a��N���iO�!F�s<��Q�= ��j�:]�zNE�����X�����G�"� ����z���9K�_8���B����I}|s�d6�M6W)�ᵗ����;�xQc=����;�+���`��ۍx�u9��HoE6�9� �r�31;?lF�)����N_�����I�4�}��_�A9tV:�ُ�-+���l��4���P�%͞���"t�_E�9YSgz�2E*�d,���u��8��3�
b�;�8r)hL��r�rלՍ��c{����k��i�>�D�Tq�i�]�����;�lm�x��P�'�3���L�j\TK������d���:h��}oj�#1&E�cc�640���큓�{���i������ps�wf�:U��*PHtR��0��R�����i�b���6�5�E��Ij��fG.��oD�p*g"�Y�95�;�M��N�b��J����q���+_(��Q���-8S�h5z=�uB�B��?�7|F�ן'��y5$�<��E(�g��޸
��=A'���;�Ƅ{ǫ��/(�9O.� �1��3���Q �nGV�pm�P)W@[���G���0</�8?���j$ӆ9Fu&�fPWDhq�[d���ib����m�zp=�`u?G��J�+]`?}���#�JCGv��"�ߓ�؋ʶL�A���mjRl��D�V�o�	 a���q�4�L��% �?cd��7Pj�Ɛc�����h�8�6����6���Q�����}�8��K�68���վ�F�T;DL����}'��o-�c|l+� ���\�
RrQ7�#�Wތ8�PF�t�ˎ��b$�	�'4,I�i"c&fƢ��KJf��i�Չ�I����KMn/
�-#�2���q�ܺ�Yg�hO����K�4)lRu�^Mt��)h�~�����-#n�#�e�IK�nW
�4�t� ��ԣB�&Mh\��S\({����o]��ʶ�B|ɍ����'
l���![��L�*e�R/�U��=�-�(��@�|�6�Z�uƒ A@T�A�$*�L����MaѲ�7��f.ŗy,��@�����.�w�o��s*���X�	�?w����G@Y\l�f9#E.�3�䑰�[ōm��s*�O��uo�	Z��(���6w���	�1п���NT��7��a�}�kB��Xb>^c�d1��f5d����U�;�F��wG�����ے֖K�s����pa!�w������͊*ͣ�iO���U1�ڊ蠠�;�����*O���h�+����G����"=�nC�����v/$́�1m��n�oKgG�FQʨo���������5��xu���銊�"��C�^.(߼N(��TQ���7s�w�I@���'>W�l��WR��#���iߪV��e��������j&��s�{ @�!��%s�̤ ��2V��~�I�tfI����V�Wǅ��S���� �0���ӧWFօW � ��''ruѳbC��8�H�77��O��o�K�=j��U��Ѝq��KҎ�����w��9�
3�5z{Xdc��,V�?\��e\K���)�GKd�V�O�&�Z�U`�j;�;-<a��I�?�N�a����at��$����Rř������Or��������գ�F����O���Eځ�P�"~�����*~�>[�/w���ZUc.h�F���(|��Z,�(��&��ұ�>��/J[tE�D�qE ���̢cM��1�[���c�2B���ϛ�;�{��`��p���5ݬ�Kezh���縋�|�Tv"ے1���� ӹn�@��jE����B����E�l�E���ʕ[��c=Mv^������z���h4`n�9��b�J�t��aGT*�����<$+�� `<Q�Ԁ]��Zi�qnإ���dD��Q�WX���`,�/�f=1�]f�ڌ�m�4�ʱ0��^V���M���I*TĊ�H�����T�=��V�)8�h�[�����b��7��Z�c�6���4���r�,K8[�-"���ŀ
��[��B�%�C~��W�&X��!_��$����*�N�3��@�/�bx5g��u٠�y��)�-Y��T�����UнuQ�n��=͐6��̍?O:$ %G�џ��� �ao�e3_!+�#����]F�Q�
��WVҍ�ēj[�/Xp���.����Y�"U팤�~;��^f��*$i*/��K�H�U9����[��3|��n+��� ^��Hb͎��Pe R]��5s(��{�@���\�*��L�UF�/�串�q�Ӕ�`�Th�I+�n�>�u�S��s�C2ϑ�n�E�p��&��F}k��G�62;�*<h�b&��	�P%�N��5m�����,��~��3�k�Oy�/���]��^쥀Dۢ5�/s�~U~6E����%9Κ?E϶j�س�n��<:���d�<>4����<����$js�����	�֬�S<����J��Yz�ŤM�:&��B�Z)K���z���ș�0���"=&H���[yƦ*{^�����5f�U�	�O�={Ӡ�5D\=�2�¼�ޓ$��d^n��4A���3m�{��p�S-m�]Ѝu��6ﴵ�1o�z�n��[O������r }��R���Ŝ�W6��IH�N܀�ʫ��4}��Io��I��`�?�X6"���}���=L|�=,s\>��R撾5-�fEӒڦ���c
�L���5!}������hs؆`gZ���Ր�y�]�f:x�n3��n��d�b���K��&��{�R���>��:���\�j���i��sH�иou�����r�b�ƾD�̞���b*��[��0��r�A�g�������5o]��
Ј��[��'9JN���#]XH(/�y�1=}	3���d��9�]��Bb���.���ӟ�Q2�"�]��c*��g�Y]K?N#Ͷ�~�h�}[i���ܞ��j;c�I��{�K-[ >/`�LP!Je-��YG\��t��aj� ��"Y�w ����uC��1�e�E�q�ZY�C�d��e�:�ޏ ��D3�h�]�F���08M��A7�����B1TB�n�7�h�ٟW�~��� ή�,�0�,ћ��������_f�b W�1�"2xZ�'=5#P�
ni��k)�,~hW�-&��
']*O�����l�b2&���h�w���i�J1��%�>;� �5x��>e��B��8y��F�}��%Q)I=���.�n�2Fd������
��g��]R�z��{���8I�k�sZʷ���'STh�}C�OK}��N��ɕ�X���Dy���@�Y���p�Ϳ��%kb����o��(���uÊ-i'�*�́��ؿ�Vm)a:KU�[����2_�:��D+	<�R�lI	_skg�P�+��7�ˠl���b&L�~��i��E�/{�Y&J8r��&�7fӻo/�tx�#�?R�]�qG,��jn���O�u���4��!&�A}��Ly�[v��'A�܊T�^�nPZ�{A�O0�'ڽ��)o� �pR+�|zJy�G�n��.�0��9�i��/��l��`Q'�w7P�+ᳰ�,s�L���&�����Ӫ�����#�Pr�8� u,&mӄ�S�hZ�jDT����%��Ei��!��l�p��
���.��CA;�^�FM�����y��B��R5�[�C�����h�5�![>p�TE��W���%���2�[�po^߯�.<vW�Ĥ9"q��a�6�c/X�*Yu�̼��
���w�S0X���OP׼��tI����g��?6�̷̙̕���@ڝ���e(�!�J7"+�U��䞠��9��5�x!��ۓ��e�`�'<��x��:j���o]�K�?1�}��qGc�r(U����;#���M�S2Q&���Q�Ů���x�ZW8U���f+�"0�S��Ʋr�5(�������݁:kZ�X�-�/�����AQ�8��'�"�ĭaD�e
��*W���JW}�Ҕ�(�,1��X.���dP���X��rg�[|�ϫ�ɵ��T��9��we�[�w!��LoI������=%�N�<��rW��~�bQ@����Fй�w�����X�x](z�RJ�щ�Ѯ���6�W±��!�\Ս��[ԉ��� /7ꎫ�S���*�G�[m��>�Bf"x1�QN0g&�oվ����/h��Đba<�7ӣ���K(�%Fm����2:7��r����>/'[rІ��w�l�]�a��{�Oe�]�*x�=�/��P��qw�{pZoL�ȝLo�A���j����B<�@�����OS����9l�¥N�
����U�\[F#���f�G�i��� (+�?�Ė��NQ���l\��B�d{��Ч����@!�[�O�Ő�WW�Ou��݊��ĻJ�q��O�LC;H������v�#D�\!�b�9l"t�������r�S�D�f�]r��Y��-g��R/��C��p�[Ò� ̢�C��w
��m��=C�y��R�������+�I��|�G.�ɵۦ��:'fzx��������)u�&��^�I�j*�%���[Qw��8��.GA��Ɍ=4ukȾ���V�!��Q((tm4�e��?M���6�>��|l� 5�([Hc�M��l����-�Ic���6�$h��5X�F^��j^����y���b�g ���Md̿A�O��|�.g��o��R��Fj�{��l��P�IZ��՞;���B�kaY��P���=�g�[*ᥳ�\�ؐ���Q��s|/�������żU����� ��:�e�xQ���㕗=��H��/b8�l�TN0$
�T�(��K<��x5/��տ��}>?�[�Ä�ex�~3֚�&���\�=���_.4��M�YW�4nR��`��J�h�xV@x�+@x��N㩉��]߶�g��T��@������]�.�U��K\�˱���f�ef1��9��ˉi5����і1{S�����w_<߱|;��d��_�7L�~MჁfr�EC����_�Sɍ_���߬���%bc�I�b�7�t�N�h~�=�}���y��Ӓc���{�7�69v��� ��e�e�����N5.4jprArS4� ����
�(r9S��^K�K8�W���p��.��
����N?=K�ՙ'C�4v,�6�ΥJ��$�H��8bL<��!�D7��ْ��]n(�>0�xK��µ�F#(�ت�F;�C�͌�jW;ԡ�WE�G]�7���f{�1�Fu�l��˙8(x�9�!C���-�l���N1�vv�N�uw�5Ys"�������$#x:`���«S��Lh�Q/�����𮁧:{Ѭ�뢞N8���E]�.W�a�:7}?'MJ��'���������#zC},ЭڌG�G��g����ܬ�'�8�/��c��f�=���I*�X�M�S��Ry6Ư��N�M!m�����%���1i��	�8�P���[�� �֭
��v�Z�T�b��#aIÃ{x�g?�܁U1nH��\#_�1�+��#��S��fd�P��E5l���-�qf�?U��4��rL���>�ش{���yz�C��6u�Z���BEP�{LݠJ��Bf�g��GXmf�Y^{;�,��Y'~��{03ZІ}���PˎP�ǧ�s��š_v#�#��Mk���АPԑE�{T��m/���^\Cq�ͅ���F��G��-ן�ŲȚ��=-6J�ErȘ��q]U��#�������M��~�
��h-4L�z�����(�%+0�('�gM ݠbL&����9G��	q�~�m�ښ�O���ޜKdD[�{��9�Vq&��;ʥz���m��/��u�%�)(��k s���DCl�Tѐ��IZ���w2x�㽏��/��N��6�M&^���4v�ig��]���4o�X"߅G����51�ކPW٧�>$b�-̙E��`:�����~�������xa�S�@�AfY�R��y�XAD�h�]���	��JS雹���1{�J۵B�F3ފ�3�ͻ�韶��Z^!�f&��Y�|9L(������p"T��r,�Dᥫ�an%�,k���)M?0`�1�>#��Z��Øak��,w�Nr��g��ǑD��*u��2�傸1����|ҏ}kB*��b%^�%�O�'��vm� }b�x�\c�6�˷+�j'���.M��O�k�ߐV����H��G)�{smҗ�꒐"I��6�H�}�`� �"���V�?S��RL=�"�h�W��.���6�'h����	�ń�M�޷ <�tBe^� ���)X�k
cxY����E���[�n����0�ܮt����\���U֦p�qx�-��}� ��@����jc����ض��W
oM���?Sitc���gt�zdB&?3���8�ɢܸbl�����'�1�Z�5�I�� RJ��A�J�"%�^�g���2�*/���/R1������ ��
��PDC5y�M9=Q{s��0�((�Ň���ђ>� �n��T�hX�n����uD��W[�FI��������h��[Ѳ�M�<��d�#@�A��D�����׿T�a��Lx]�'�'�ʃ�[wY�DmhF[��%��O��0�5j�]�Z�y�Y(��Ҥ2���<���Ed���>��k�;�g�l���F{�B{���A�7�'ǻ�w�oE�1���%�ז��e��T�C$�RN���,3v67�D��*'�gt����S/�g&&�����!��]E�Fi("�jL�'���%�ƽ�ճbI�%!Xy�2K1�1���F�yy*ٙٞ����������|�de99n���[m*��#!j,���Y��aPHԝx��Yпw�V>c�-�)MVq���'��y���i5T��RK�|/P�i2{����Ŝ&�J�f���.��;�Θ����9jKF��f�5�Q�|��G���'�̈���Ѳ�J��*�K<w�$պ�n�-h�S��eR��Lz�s08�(e`z7�a+F'H�'/d��UQ���p�]Bٍ��x}�5�[����T��jM|ٖy]��)�6�+�n�����32�d�@�j����l�v�
����ˊ�ㆮ�r ؘ{*����d��(�@�N��Z�ޓ��ǁ#��z$�	DW���	Cn�ů�V������{P&a4���/k5X�c��}t�~Q��D+�y�;`hG��`B\
�I����	�w�$�2)}��o�9mKO��*�D�"fOp�P��9��~��b�K��~s�)ňwu�g5G�>ek�Růn�u�6�?��\�\��>!�|ַ�ƿ�Lk�vN�_����5�q��I19o8��Jte ȋ�MG�2&�o�J_�Ċ��m�I�&W��g<��_�[�k��3&7׌�
�L k��9�,X�,q,a��#ڱ=�u�2����_T�mN�~��t;c"y�Zs8�˪m�O)n�_��Ͽ�V�WQ�\Q�$�E!3�40�*HC�j�J���t�����q{�~�{�n�xCc�iӥ�;��2]@	U���ϲ�L7ƕ����'�@�X�rU�v�l
#�����Y��8e\�o��G1����?�����{�� ���7v�pY�{�%���_4_0#��h�lm7�Y8 �[6�(�K�OT��T�3@d4�����}�}J��<���r�ԉ	.�t6�2;c�� l����z�@��A}�GF����RH�\�V��f�i��)!�ɂmF�����wO��}*"^2␱�w��{�1��B"�]2�ώ����ة��B!�)�rcΓ�ǅ}�EL�ڳoS��ih�gd�#l"�R[t���Nv	'#q��?�D�ynv����@�-;�d�n�vd8�iH��5<���G��L%h�����{�f��|~�s>�|Ғ>��cm�lgGdr'd����#��y+"��}��Ų*Uy�s���!�)�z]� ��d����������R�a1)/��=7#��`�SI�oH[� L���7B��L�T���Ư� �wI����uM�#oP7�:�j�w��hĦfǜ[����ݽ� �&7FưQv'����#��iPN ػ�=��c�x*<��ɡ/�)�k�����aaݳ$�P��-0�Xs������ς]di����:]� ���z����SVH��8�?�.!p�
��{� f�Ļ0H"K>䣂�,�켩S���j'̎(�z� �������i��3�W3�.�h��L��Y�Oj���5!|���9	C�W�O��VZ-'
���4�J�����v��є'�׭^���`�8��BG
�ܸg��_����*b��5j=�,S#�2:����+he�ډ(��rE��d���|M�-ZBq�=5տ�TCYf�*�k%.�ɾ���|Y4��`u�o���H~C!Ϲи�!�j-�.u�>�&��t>�C�$��d߬�C���J�}�6gC����]��Ϧk�zUk-���x/i!���4�2��oo��U�5�*�QŸ�21�xLe�I:���8���M��X�.YMp(��h��[eb'��_��/�A��^����0�G`��1`�"MwP��vƩ��yW�n���%��H�@��+����!�.�v��s�X� er���"!?�ߓ�jl���5r�6�U�1%ݗ.�fɺ ��LJM��2��7���Ϧ3B��[��W���(�"�o�瞖sb�x#]����Td�Q���L���:��������fa�P�O�)�sZ�͆{�.(���d���a�ꌑm��s*^>p��^A\��1=Q����'�*soBrW���EڳWeJ�ڦ�D	 ���{1E�Q��/ �L���9����6���Y[���'�WҜ[��mcX׉MnǨ:&&�F4w�E�"�Ak��ζ�.nf�P��sA�Z�D��'2�G�F<[N�
�����|OD������p2�(�j�����#2H���?t�Q������'m���'�B蚛���u
jǅ��*5��T}�FFG>���*�JG��z�q�����kM��y��6=��'�3G�톶�&��~���$�W�j��7�
�*�ZG���4d�9�@��U����.s )M�V�9�WRL��ϟ8Q*�=T��*� ��
ԑ
+lRX���7���A+����u��m�L��	��m�h<#��6S ���ƂcD;к�ts�yU��3�;�ݘ�n���y��! ��ߐ~"��-m�X�hۙz;lML���9�f-lH�8��g��x�߷8�J^1)��X�t��C�z��±%��uԍ��t{%��O�*�hK�RϘ�E
a,�S�]��Gz�
<(" >�!�;�Z��lN
!;���TO�>R��T��N����y����sF���&x9�7��C�R6�F�vw��Up��Wg���~0�=�'(�n �<���}\g�^������{��~Q�@]����%k�Gb~����ep�(��e%ɇ����.�hb��ͳ�D�bc�y5��E��P�.�~Ssؔl��3a�X�^!o*x�M���!��.�����C�D3�p�u�ֆ�:�i�D�4l��e*�� ��+_S����=���LZ�������j����#i�Q���s�#Zaф�����&�"��y�ɪ���P��7��Ι��Q�C�˺��maNv�v�;�}ȫ�m��I�)������)~4�G���v��e�|p1V�Ӟ%b����6�Ԙ�4���v��j �E��􂝄�Q	�?��v�9 #x��=(�z3��#�Rr�D��u)����8�X�=�ri7��0Vݻ�LF�]v��A��_��j�>`�l@)��3���ي���hі{%�&�����\�`>	���F����.�OI�G�D,Ξց雄�R�,��x��Y��u�S�p��%�T|���c՚c�i?�?Q6��0�c��0���`���	����@'�(��m2�1
�7��P7X�{��*Tu%��#5K*?�����:� L��������X��HNlPΏ8"��V�=�/�g���H���^1
�a�i���RE�9�x���y��C�r���B��`?�
�%�uJLG�>O$Bړ�˒�7��l����� ��X�E���T(�O��J�Hfl�p-�F_m�0_e�{��9�O�$KǼ��R�ߐ�Z�N=*ݟ���1R��@����`�����(_�)�`\����d�r�c������-��H�� �#��/��lH����fL\Q@W�,쐐��G�����Q�������K'pC'Y�Ю�)���|G����~xS����L�@!r���e=��s���RgUl�pnغ&���Uy3AP*ܪ�����{�ى[V}p��=A��r֘'7:�;΀��3~�=��A%U����g@�X��4	 �Hs��ECY��{�)�=�\�|���[ے:��}�yV�t�4�ё���h�y�޷#��˔�hf܊�M��Z���|������վS��-ߴa����A���V�z�����]옳G-�j�܂�ؐ�(~�DY-����o�_P(�>��+ބ6JK��fÇr��J�n"p�T�y��2]%H����t�7�L���g,�D���XS�A	�2�@x�f5��ƳF��`c+(_x��Hg���ruO�i�

�jz��
B=^6���(�8��"�����C��-�Mٌ~�v�ܯ+;MF#�?c헔{OI�:dY�t�?�w�w����8�@4����: ���:m��o�`��y� *�AD��r�Z"P��	Z�o��	�j�eg'd[�+�.��z�I�V��ͭ]ߺU�/�
���e[w~��������
��qtr�p��G�p��a�7��!�v�jok&w����7�2��l�%���#�=|�[s�eT "�� �Y��o�f#��9Ow�ѓ㸔j�>���9�ƕeJ�K~j�b�"�	J�ߕ���ld�Qv�������vX�M�{9�s�/�-y��"�e���Rz��j����H�@��(]�����Ɂ�!�N?^oj�I)����A�2���wU�晟�5����=���:byB�Z!Ma'zg��X�F���Ϟ�dF;;9M��{Ѓ�ʦ{@1ĝ��X.����L����3v�z*!����p�V� �5�IHK�W�8H���-=BvӁ��U����0 ��N��^�lZ�$,s�e�8Pr��Kξ��t��Y�g^U������s�<JѴ�P4�i�&Wc�\���ȥ�-`^Z�덐�`� P�K�G�[o�@�^0���Z�d���1l�+�Z�! �}U��̕����0��q̑Jn�t$'6�rr&RrQM�/�"��@��5��x��Jf�ina0��Qy� �� ÷��[�\g(��%:�� ��I`�=z��kxYaѫd�~J�g��f��<ߐ}��+��e:��y��� 2��2sK?V�$�br�|�#����Ω�k�j��r����53	|P�ڋvw��� ����������7R�>���lfQ�Y�RWr��u��A4k������SѢ�J����ᜏ�]������<��4B[oJ~�=���roA����</��J�g�{�T�v�>���6�I5v���6w*�e
��$[�U|E�U;��>��ŋ� |kTM.��*�E�����$X���ED����x�Z��0}w��&�j0+�0y08@Ŗ�p�L�GQ����� 3�
���	��Ŏm����f��*���>��#�s�c_L�<��]���]|��� �;ثa@.F�¬c�Ji�&�����Ƌ����:~[T��[����j��q�k~�,�ICvw:�'z1�
��d�̺�i�����5�Y�F3�ey�QA>Č�7�4�nh5h>Ej��� ����+�� N/��_@ظs�/����&�Iۛ�Q����P\c8����f m�/���@�X��o>hz�~j�'Z	��ک�q-��	j��ȍ�Y��}�����s�$��J��u}UCAt���P����~5�+8Ծ�)��֣
���>=�^5o��g/53�P�B��zv�)�K	�D�F'm�{5@�R��1��Z��bd�������B!cǏ��wɰkj{�\o*��}n�����hfp��) ���@	�&m�f�6k͢.���ROl���Ξ�s@iհ��0k��^&N(ӟ[�HFr�80$��P��@��:K:�[����Ґd�jO̿������e���-��	U<�ƨ54��!cc�� �a�|ڔ�'Q~�q6���Y��-ĲQr���Y�J�KIF?="<҄������9��P*��ȕ�ܲ%jMB�ů�ku�Y��E����LGK���q�(o^Y�\O����ڪS*jCG	Z����W -��������z��k��#h�W�>$>��F��`��*�I)b�W����p?��Ӎ��E� %@w�bg�u�O�u���X� �8@�Ɩž��e�i��x=�D���[���(���-�S�����]	�}�݁`δ�!��J���̛�}/�FA*�U��2ي/��7���Nk��l�~��	�K�e"�_C�D� 9����/��j���r�t�d�M�"�h���҈�D�/�w�S�	���M�Bv��˞��Z l�̒a<G��HhK�l3�Ω�Ώ&��P�B��J�	�[@r q�YA���;��ZWQ��݇�i��*5
P*�"ΰ/I��,qJ�� �0��=J�?��Ɍag�`�r�n��>s��$��	�C��W%B*�Yd��>��晇�i�v��@����)�p��%]r�>����D;�:����R�NqjQ;s����$y�\$�,�"F�D5��$?�LƔ��'�MT���]�_@�[ɔ#��>��~���
�P/Ө�)SŪt�iwUr�:��;�ŵ&�o�Z��GO�ƶT1����l!8�c1�jQ��~�-�ګ��4�9���P��&Qs�@�#f��'8V�Z��l�����/ٚT<	�[��B��=XϯY�9������u�\^~Ю��{ZpfW�A�Zt��S� '4�L?���/	AL0����6����6���k�M�{����B��u���[5EH���3�������91�&;�|����������'<�*=-��J 	������LM{Y��jά�vb:��.����2W9�*挞P��)I&�C���˭&�uՃ�ɦ���%K�.�5��gd�~��"��{7'u�X���-�K��1��#���P>�Ĥ��)��ng(�G�Ǔ�29����l{b]�~��b9�ɣ:q1V;���XGE��"�}B�&�w!`�����b,g��3$aîq���*����j��W�M�/ȳ�g?ia�D �����gz��y^k�v�Ǽ�A������"��[�FG�,�U	\U��Am�:kl��7àa�m�%:hU�&�r�R��i���Gri����u�c�q��rŝ(t���2�#X#Ֆ�An��IC`��q��t�Qh�*Cy5��5�j���߮wL�=���|``�'3� )B�v;��֕H��&��\2Xİ���7$A���ya�z��N�6�/��9rg���|bL�SI���-ң$�Kʧ�idq1���P�ރ��0�d���j�q�VA?�Q�Pl5�dW�77�=�H)yݷ����6�b(�оO�Hh�����Nų0��0���I�����5i'���(d�Ε��0zF�Y'X��G0t�eVj)�z8�s�����LMa�I�[����m.��! �p{�#,��]
��	�_�N��7����)!Lk�Au�Sվ�>.��,)X���*?m.������6�Z����� "3kƄ,�W��X�~a�)��]�Qj���i�?��!���u'��0�N]���y8RBZ�,.$G�c�>�������_R6�gO�=�n�p������;e\[��y���Mٌ?e������p^֠7��.�Q��C�/�Ù>�|Y�Q�����2zB�l�n�����;[��y��v2� �<L3N=45���ܰk��.᫨ɔ C2��NEz�-v����->�8�ҕy�X�=��q.��d%)��;�:�V�KY|8��
�.��J,?��
���a�$|:�ut�!I��ލ�bB��Oxߒ/�L�7���J�������g�*�
u�*��ֲ��4F�Q���s��t&�/���*�w�vm�_�~�f&��o)umwL��~2/G^�n͎� ����I���RW*ʳ�o���CK3�KH����e9W��S�@6D5�^x~��J��)o�b�"���b�d��|\�K��5\{ĭ��,�A�C#j��]<1�/�8 ]CU��]��Q=����s��5��Bs�������!��q��n�6:���wC�@��F�\U��0?J�WR+2��l��rt�dl�ԟJr^��y%z�횕/\Z24��}�*�^X%˪�[�m-�m���'���������3�g���I��k;�Z@�j�h-{����*g�w	����v@��43i����h�v����>��9�v���c�(yNfqE;�(���ϲ�R�sMr�k)x���~r:��ֳ;�w@P�a�	�`�s�+���"���O�4$w����D���';>Xc�����~*	����┎����D�<ZpxE�7#Q� �[M/a�u�r�y�dD�����׮P��l�Y�p0����M�Ca!���{a�S$..9hv�i�#�����B��m��׈����,�5eS,=���]�~X+pE�9L��ܡS����k'��D'X�O��D���3s��u<�u�2K���my��q�6kk�����6�Q� �t�T���=c�����j�w:+��JD���͗c��b}�Ǧ��<w����m��u�s.r ��m#��N^1ZPG���G�8�nСV���Áᴞ� X>�C����f�ّFBW;�@n^1�n3v 9��"�o��^D3Qb�Bĕ��4��K�-�'�Ԇ]�T[�+�J�IS�j۪����C8������u��Ǐt�]�{1��0Y��V�㛰N��t#S
зX�,��&Af�#�B��ה]Ѭ�&]�uut��d�:�z�x�;�-�R�}{��΁_��h�f\d��7�.pS$ΙB��^���S��{��V�aS�6,
bt�ؙe5*�@FLz����.%�	���D�}�SȻ1o)�!N�:�����
#�}�!�
�� ���:mv�6o�P��;f�*��O5�[G5u�OFI��_��K��W�ڟTDМ2��_�2�.�Dh��5�����:�)cKm���αr��v/0P�䐷Y`B�%3w����%K��LV����>�����X�"���H-�g	�Z�h��n�<&V���Y�4מ�& �BU�Gd�SW�B���|~{����K����*���.H�@��IVXd|c˷x�<:喝Ŗ
�"��hq�t�j�!F_ȿ�ެic"��p�iT��֙d*Gȁ������4�"(�p��*��{���}l�;1g���+
�pvw��ᱜ�Д�X]Z���92k�n�K�1�&�ѷ2Fc���e@�sN���꒿Z����g�������(���?l�T�_2&1O�re�i:_��a[�ɐ�\�K[�$�P`![j�˪�\-4x�R#��G�	#���_سg�r�[V,��m�����x�<zW�Υs�Yy�E"������!@�	�;�������Q�l�x4�
���f{L��h�,��:���׶{1� ���
pX�9S��`����L��|Yo%�%Bɍ��Tс�9�����xε,�h/ԛ��\��;�m6���v��=h�n�]`4��ڗ�&��K٤ ��
m����o���K�7����0x�[���x�A6W�IW9�.~�nV�!Q;YȐD� ���/{�p��S��7�n�8�E���Vp�&]�>�����g�h��R}��Ӑ�s��}�7CGㄪ�F��>��Y����[��
,�d ?6p���%�n�7�� P�K�Pm�X��+���~�H�L$�a�*����nM7�C�$t� v�
@Iq��Eܢ ֱ�y22�H�~�l2lZ�!�\�k���w ���;�������e��V��owtk���I<��h2�_ZEBt�%Q������\����.��PSd�b�۔�d���G�L��F0�'i�}h/�C�o�{�2LF� V�h�0�N�pF���Y�T^B��ۄ7�
�o����Sh�ڌ�� �D�s�W��	jF��@���1��E�����Ἴ�>�'������T��9P+FHn�P�-i��U�Bو�����)�Oڲ �����Z�o�|�K�kS�2���q	���;�b� �]��B��b4��U�(HyR.��(�`�ab�ՠ�<���R<�*iՂ�\� ֭�^�'&%C|�� \���1�}���'�A�zK�:p�'N�O9�40����5y��y�G�1ĭ��iׄ��f͝@Ed�r^2I�|�Õ�����ۭ�";�
���\uD�?�g�)ԫ��� ���T[�P3C����T�ꁭ������}i�?L k��f$�w���I �򋝩���I��먼[/*��

�/��w団�@�e��r��2��3�݆6�Uq���&� �����t�����mвt<:��J�,�)7����A{�����|��s[�)0��o�w����ͯ����EV�n�E��%OK�[�������>,i�1���ri�>��} )_�2I٪d/�!޹�RK�m��4-A(���9�[��%"!�to���C������F�:�)]�Sӟ	�oV�(F��+`'��-ltJXTP�Ա��`?�_m�A�tF�hV�P�.΄���<
A�/���?�Kfw����� �md�^�����!�j��2�a�	6ļA8"��և0V.�p܎H8��6I�p9��xI����4~s<�㈔�-3�6�����_� �i4���?Q��voh}/5���ɽۿI���26=��)�j�����K��j���(������^2�'|݈HJ���ۯ"�b�8A��.ȉ��@g��M�� �[G��nHՁv�T�#�ؖ�����^��{��9�ɐ��_��TJ�F:��3��'ČS�L�^�nm�1Z�����-�"F)��Ʉ] ��D�N�f�Kq�iP8�ꮑl̛|�/��a��"�vE*�Rt�m�ڛv����;�2dS�ҙ�N����ƛ�P�nE4�ӜJ�f�9�W�ݵwSi�X�����bjh�x���Meղk���J���t�#R�.��(zQ8� �J"e)v��O(��g�9/�7�=4�0��Bk��F"o�;�]!�#�P���
#T�`z1��'��|�%�t�́��1�8�zf�f�t�����ّ��	r��"����r/ޛ�]R��ɪ�y}UZ@mF4�r��B�sg�q�yzSJ�-�e5ؾl�7�{X�:������&)N���/<���Ktx�Ļׯʺ�1��
cÖc�� A�%��������L��#�)�d�]jOZ3��>r�ȘI�V<�q$21��[�z�ґ!�sϜei�"�d���2��B�,����YB���2�A�������}�>��!d����U�ޏ�~�2El���cG�����Hs�2���p!X�������c"9x��_Cɯ�y��-cg��?�$�5o5�A��I��-xߗ7kJ��+hS�}I9;j����zlFk��q�nP�[�g����|!#����⹰Z�&0�����!)� �������G�n��S�{��x���Ć�(z�	�}���
�Nww����:�wj"����L)[�#8����>I�!Wi�A2O@(͙�Re9ڼgz�M��w;kG��ǻ-������39K'�U͖A*HJs !%z+���Tx��%.h��mL��$����0��k�_<��I��A*��^���<:�u��4�O���wk���c���d�l�
�q�FZrlY�2SrK֋���fY-ja����ZUqt�D���P&Ya�J�I��ÅxX���Z�^�r�L����<m��a�y��%���:O~¾s�)t�B	��exI��ue���1Q4^͵fY�tj�Y|sfc?��2��>Xq790�^٘��t���-xY�%z�D���Y�k��`�:+~�>�ӽ3�+����%�?�����T��Ⴟ����ni|i���t9u������9��I�o�x�O���K�_t����U9���7L��0�,�8IcZO��#�ى'=��(p�q_�q��+~�[��l�������������#�À�X�F�!q��sQ����Ǝ����yL Rǭp0Sf�튽�@�\�(�;w�����{d2��Z��0��l]g��;�,�pg�#���s���z[^�)-/�-5d���.ȴ��2?�ip:���$�!�������ϓ�	6�����!��\���{Q���ǧ�-\���?,T#�YM�V�,ݧ��3N��˻����0�;���5���Ho،_T�����e��M�wL�̴1	o!����9
��aP0���!�>�i��� ���P[�vF�*��A&6�� ��́�:L� _9�Y�A�W)k!�AS�v��R�3�p�����: ~ԣ1>J�@�yx��BGЖg7|�9��ۣ>UP1j�*D�g2u��"r�Igx�ŏ�Ħ���o�T��r� Sr�r�xO	�h���\,���@����K4wFU�=�ey'��Y������s��R�~�R7�1ҏͫ�~���R<'�9�螊#�l��vAvz���coO�8�[��LvӐk�)�0�oD��]f1�V�?%�UvuJ�.�YZe��60p���H
�$��ӵ
�ǔ���Wir
qW�I<�c��`�i��n�w����&B>�X�woF��)��$m�S��Ĵ�(����1��h�E�-�/g.��!b��E6-�=Н[�G��J1I�O'5�.� M3vS���]�ߧG�_��f��^ZHՏ�pD=���κ�ݪJv���VR�	F��s��U��o�oa������K���]G���d��܉ӑk=L�0�+�*��'�E����|��M�Zӳ�����{�ɻ�J]d� �.��@o?�e0˚�����P��O$��7?�����h��� ����PtCD�L�ѬJ���e"��N$�����V��O����|��Hm�.F�t�X3k\�vg'-GS|��1��ٳ�Ќ�F
��M��:�!i��3�C�����tMV����2P���U@S�hce̤��ѽ���2(���6w�5G
]@���_�*b�D͢�͢���]*�ɔ0��X�7�(ԁ�0M𦾍&���P����%�E� �+�i�+�?׽�����w�o���y��B覈��P����c�6�J+��b=v�3����*0v��c?j�x��:���:�~����B#�bpj�9�hq�HJ�lB�����1�tUU�#���N����u�#����&1�\��MW�g��4�	����X��wMq���F���Y`���d3X����r:I�%��ê)��� �����6�e6x��QWWi}����+��f4��%e}���U' ���!�Zמ�#��a^���ӳ���;�Wm��~/�����;������EI ||�����L}�"��6k���Q\ ���m7�5)��뫐?����B�Z�4P?V}`���_E�ҟ%�N�N'���x@=K1DW~�wB|Q�U��D������wfmbJ �G��ZT��p+��V0H�[�V�����ݻ��a��wIo���xB�d�bU	������>�\�_3~�ܺ�c���Ȱ#!�0{��8�o;-�e����`΀�߸L��'%}1�r�C{+NEƿ�KMo�̰���]锉v�1{�-H:.��ᒓ�
3��j{Ow�U�1���k���|����;���e_/�����?m���(��oNw�`�ۥǐ�/�@��j.W �0ђ�M�f���^r��}�76�zq��4k�p���7B���c���c��Eh:J�L1�	�'�wh�2=�E��;�1���6������U��#��w� �@���ҍ>u��־���][�x�Q�>2����q���q��Ap�ή��YW9�,����y�=� �	��!;H���yw�&t���t6���� ���qb����i��ZW��5+xK���f�4��{�͚Ѩ���B����x%e�븝��}�������EyK2�p�>xb�/i�l_���Y��V{\�*���,�!G唓�j��Z��=��<��$ơ��տq�[���㺸� !�P���
9���I���
��F"�����9X)�a��,oO0�`����h��o�] �rr���	�2��K�0m:mP-�I���+sC=26���� L]�O�#�XY��❏W"�7"���v�f�e���is^�T�0�Q���9��~���*���?�)�D�d�Z��{���gH7�u]��M��L��
���=�-x|$*�e�.��3�����@NYA"r�����+�s�;f�R�I��.f����D����Z�����'�E�3In,X���`^�i�~�(��c��y��c�&lC��f�F�Y�t��K�DtR2����P���צ8`�l!��L-�k�2�>gMXF��z�G��z��is�3�(�y�Kl���̹��4̆훉Uj/B�؈N��'�s�|ǂŐ�IK+�Ld� �~Z�,b����	�t%,b+#{
�._z�s?�MKĺ�A:�SFq0�^"���t��%�S������.�
8H,��-��mzk���U/�����}7wV>��O�P�+X��oSV�}kT�Ii��F�0_����T��
\8�ŭ��zO뿳���+����N.
�,��߱������+��+�fls����Wx�*1SA��.ŝŮ�� �֎I[d�ܕ@A������M5,n=������OWM��r.:<��ׄc�]�D�j&�xm�6z�6B[���H^
6���4U�.�n���O�
��Jkȶ�	N���3*lA��J��xo�?ă}I�sX;iӛ��r.���gç"��g�|e�.-�#Em�/�6��c��ݜw�!BKZ�\��@�i ���cF-Mם������an���J�y���c=��`Dl�itc��_���5����~����Qc�����@��.T�d �)�29e`ޯۿ��ك��G���۸|5����ئ^��g�lJn,��yY�4sU�Oc�x#t�d��2�d�tw��S�:k�
���}5nH����tx�c���(	�zn�����e���y��#�A��C(�M�ϰ>�҂,�/+�+�44�I������LbƘ�0��S�+]��D���o���ô7�Aמ�6�h�s�����Bh�9����]3�2Txf&6�����6^��FH*�P;'��z8����1P��ѹ��m�o�1^���ٿ�[��0w����c�Da�5��<���tqw33Jݩ�kd�ˁ���t�єuF���ߕs�9a��m���'E���E��)�c�&��h�yF�|��b�&�YSJ�<g~��� A�F�&���%$uU� �^���&���둴j�,���4ˀeLiX �A�Z�ԇ�`�#���M��q:`+��	�;���Llu�%v^�z�
�Oq��"�j�)���jC���f��Iw_�khc��p��]�Qa~ �3���S�q�%�:#Ԗ���ؔ���;������˨b`���|���7�i38���j
��(����W�&��j�.�)B�v���/m�%���%]DAQ�Q+*�^��5AQ��+�+qT��xD�Q�z�Fh:Rv%�9���$5�FQ�Z4�մ�;EA��CY����ԣ؏�`��_�a�9�}���x�0�u����e6s��Tt?1^Ь�L3�K��z{� I��ק�MM��w)XI	v=
݌,����P�k��-��r��@�z�j�856@�9�Ky��W|+z�&�k�3��߮�����+���a4�"%i}�9�M"���+-��Ӭ��+�#��G�R��?�^km�.l��Y�JS~�y!*{v�����O<J
,M���j�+~�^�D�X�Y���4{f��O8�)Kz��Q�/�
�1���2-U2|�>D3ҏ�"'
��5�?�~.\\�	pwS��C��Vʟ4�"lOc)l±��WT<�`��L���d���2���]x4�N�ps��C�#�����u�JC�(��{
K����32���.��7b�^�;�}~���jJ��I	lc$�S|�Y
���!��+n����c۾���M�	&�~�e�Kn�mNB.%[ȷB��#v7�*Z����K�+�~�(��Rh��QI1R�#���{�M@�����eNo������9n�D�%�D�*� r��d�kH�����s�I�♕O|��p��c �r��e(k��*�����gd��g�j����RS�e5\&�M�d�2>G��O��8���m��ve�Xf�U���Ԑ�R�fV{��O`2�qdh>�6�֝�-[������ݟ��%�Nt�݁�a�$f��0�D>���׭�"q�]������nX�� ���Bpg-t���d��.ǅ�܆f[��:�Ѕ�j6�J�3'cT�>�bh0 ��Av��bʼo��8g'9ux@��N�<#��W�\9�U�U�L �jl��y��y�:����oU>@���N��u�d�Z���2I�~P����Y�R�s�P����A:�� ��U����W��n�l!��X��6mr��
q�m��%W (	�`fA������C�2yEM���:K�a��g��˚��}=u�F�>J��ZkV������:p�t�6 ���z�7��٨g�VK����q+v͜�R����s��J�#�U���Uo��.\1K��3���w�!�ӊҢ�}�d�2/�4�zrb���(�PW�C���&�I��褃�k���Bg�2I1�=���[�JTU�ɥ^P�;����]�
]�l�t�}�׺�vE��Ѥ2:�|�T��vHz �����B~{��[B_e.Y���������h7�O�9m���&`t9��_�>=��4�0�g��N�Sf�j8�X(f�f�s�'}o��?�|�5���dAvj3Č_W�'M��J��:*J�\����ޘ[�ׄ9��{�&K@�>WB�8�fS���/�7�
�w�?;���+A�0����"�� �C�P�f.��K5E�����tϏ��x~wIL�u��[��Q�[��q�f�e��,�)�&�.��h�5v�-��E������ݟ$�|�Az4кbx(?�!�0K��##�����9qo~o& �J�H��]S��鄙+w��o.�G@�$'3E�X���pn3L��M�7�:&&P�#�~F�����`X�m��z�z3�z��\��@Z�Ϳ�"y�$���l��ԇ�;�i��j�)���x���$��]$�,�ܲ`��Pt)ZH��P���8)3)�/a�c��d��}7��T=U�VEsؾ�N���*�����d�`����f�1m=mOU*� ifҊ���C4H����?S�N�flb�
�@s�c{�u"L���ǔbo��#��l���+�tP�n�&'�þL|���.�2m��c�ߥ�Q<�V�2D�d�{7�9��E9��$S	l��cm�!r��};����z��i�D򝲡�<�N��B��ː��&,������ʰي�\Χ��_w�(T)&���G�X�G>�Al�c��i2�P�N��#�F���xz6�B�򏄀��j5�V��51-� � M����Z��[�9���<������qC��ScY�ξ[ioG#�@rb��o�>��bʊf{����7�Q	:JtK�z{�F�nwe�q�}q��*_I��{���}K�9.�̱�1�����r��6�H@�U���\�J��
�?�L?�^RӴ�6��v6�͜��à�5��z�.�W��XߢQ�7�.?��P+'�|�<����a,���|�[cY0�Qm�_m�ˠBD�w�` ���	+�#w"N¨�s�m@������9�S��L}�7�#;�k��a[��ؐc�V�#[�R{E���V/���Ǿ��JK�]������P�t�iTkh-7�;�	"P�À�I��]~v��D{Z=��~��V���~謚��.�
<���'=�a� ���,�4䷔�o��جg��ci��9���I�������Uj��"�Z�/,�����͆s���p�t����c����I�#�1[�i���y|�#pP]iS�v6_p���\/[}V����?m�	b��Ś_�'C���qg���1p���BiXq�'���N�V�0L֩���F��		Ѥ����,�wlP�ۭ�ha*�W
�0�(�Ӑ��t^����R����m��k�&����� {�ԤCbGž�[u�7)�S7Y���Q[�u�Oy�_}��B��b12G<����`P�	��BtTbj}k���!��~�hF�X��^x���\-W=��X�����������gh��
��t�Q�&4��%;K�!�.�)�@���1�F	3�]����7����r�fH�$lbK�Ͷ�{ʝ�}������Ўy����]��#�$����=�b�ˈ�*D��]KS�h�*��5Z��I���稫�K����_�f��$:�{��rM4�jt/"���ԧq���2�Q��X�J�Z��9^�aRc#k���2;�E5ѕg}���<W/ke�o�K*-p���G
ؗ=vh	�/���A1��e�At���`��x�7<	*@ �=�S�����,+"��r��n�.1�zP��s�<��b ��N(�g%��+��=��;�� %�8��=�O�
�������H��%��|I�rN��3�������ZEw��wڵ\~tE[�ً��N��1dj�ma���Y4-1�u�G[�����*���@7�H*���9X��;zA��+�M��\���z�V����)nuU�l�L�+U�S�WՊ"W˻ɾW��	��X�Ddj4���\mˮ�m�^m�SV���u����E9� ���.�����w���6� ^2�f�,�g�Y���-d���0�L��yU"̩41RMb�[r�FeD���᯵1�Xj3$x�W�/�d^[��̫�9=��VV�;�jc�b����Xу���?l���Z#'%NP�e�fa�����1���Il������Jp��|7K�7u�:����HOiJ;<����:��K(!ܩ�g���*6��>�
&�႑�����l���dw����|MC��Z��G�k�C,[Ir�	�Q��,oӃi��(f�6_����z�>���@�C���č������ts�����V��#��U@M)J����J�� d(�'
�g�&�V,h�d�៩�H�'�lbU���u�:�Ӊ.~�J�4N��qS.�?��_k�n����b��EQ
}��y�̙�H�'����8�5�f����q��Y�\�V�m�碠)�
ب�iu�b+��x����ԓ�h�vp� �0FJv�6*���B�P�9��(ߝ#Z�>T?]����1��:�_��7����E�u�Ð���(�ߩ!��&����-[h�e}�����t(�����Q���"�����>����\��L~ì2OX�Q�j���M�L�HI�� ��r"�a;����%R���rK���2=fH5�cp�09��Ne��#��M�Q�nʞ��%JI��`g9'?��p�L�B�]sx�I@��Ej~w��l"����̄���^FEw�c�[���R#���R��1rm�2gj�hh�ڗG�@���u�ؐg���Fn�tae��q)W6��<Ec/-�<���e���qHC eW"W&
(�2������EH�R������d>a!W�\�vr����q��?V����5(���]��H2]&ӑ�(��ڴ+����.�E��#Ny9��h� K
����f��j��U���hs�񏲖x@`q�,�I��k���S6k�%��
<��(,�í-�|�5o)�$Ѿ����w�����ݤ�� \/5J�M(�v���Z�J����y9��c�O��Id��Y9#���z��T9�����d]st��L6�n1v!�q��3���6n���+�K�Ĩ�g���k�[j������.�z��]�w͎̃>GO<0���7��!#(��XY�����e��bЉf_�j��U���c?Rj��%uaT���&*"uz_J�7d���=�<
���+GԼ��ؚ}Ǫ�-�"`x`�7�{�Bc��&���T,����Z�Rii��o�F:��=�a!��3mO"i� �^�W�J,$���[�L�L��\�[�TT�,�Z�n^l<	��Xe��i��Z��p4QFD&'��"Q-v+��4X(d��L}�#�jNz���1(ѣ�)p8��!���F�̮r��'b`Nb�ț����6�O�#�ܜ�j5J;���E�&-d��	��h���]#h�K����,؝_����j�oc�MS�����ex0<O5a�Z(Vm��A)&E�c��{^�d�^�wk���?��?�?�7����-�;�b3����}C���$=��`��,`�*+ߊ6E���jN��(��{��v^�˃�U��!���z�����k�0���&�VbfςZ��qE�A������<w�����/~��Cꛚ�r��L��K��>�W#0 :��c��~�/����>�<0kHy4��SoD�\`���*�I"%�\F}�޿�iI6�G�A2�������m�(�#��O���0F�6�M��'I�X?}�4D|�����RK�n�ַ�V�6\�������gR��p����Y%�W�5]������N�z����lT��wΈ��RoeI�.���H�Ż��7�(������P$V��(�����Zo�U�=��l��ߔu�s���6�ik�TS-����t�(� MI#h/��X�j3�����e%�����~��>[��	���NY�ݟFH.'$�߸"�����#�1e��P�;�{�ȹ���Ң����(��R����	Q��[�.�;�R�C�$y�c ��4i�k�\��� x�,�T[��
`xm)t�￮��})b�̍�y
���)V������@y@�ux<�O�l����{e�ᆴ�� #����i�X�B�}C+�z�'I:���e�@�P�Kt�����=-��%D�r�6�`��$�?'le M�mL��ϰ3Z�[�M�@*W'U��>8Y��)�q�� <S:�(�'P�f"�F D�$���s�?�7Lh%@�-�1 K-ɜjg��s�忡�����W���U��<�����1�W>0]ygp�
�����!4�[8etЦr�ǝ��xI~_C�˶J�^
��~��E���	��Z���J�c���i:�f�nR���\�����*�.lʃ{;�� ��y��?Xl	�j0���o��Not{�'����跂O͝��iJ���*?I�#��S(e7/����a>;��B3MÅ��N���	�2sC�Qa��A�K���Rl��m1�,X�4Q�=�Qr�����@�Py+�G�*�r*��v��L���ɼ�*�$�����"�c%�N����yY&�MZ��Ȅk�WSa!M�p2�v17���?����ʗ����n"+�����\	{n�J ��<�eظ#��_q)�÷ϙ	��1�a��`�
�~b�G甌�ߋf�y�ҁi��P&�U�H�%�����ѷ�!�2Y��+��,�I@��w��v���?O�2):�I�;	R��K_�i�zI���n҅V��[SǶ�T������j��[,Q��B?����#�B��V�����mh���;��4[]?�Q���}� ?�S���mm���S�<���J��6\���Β;2]aF6��ʯ����uw���ƬOG[}�Z�ܸ�-�+��8���I�_�z���Bί'k\Α�Ϣ��-ɵ_K�}O#�o���N#��B�z/��F*}M��"�xF��*��#��U��)ϯs�ݪ��0�iV�hQ����f0)T������O ���PҠ��Ƽ�>�M���R��{D tk)7p7�;�G�MP�0���q��36�)@v9�Fl�W��<�?�P$6�z4�,/y�����Ob%�iK�7��� A3���������i�)t��D5�Z����1҈��t�{b�����E���M]�����L38Z�N�A�|���I��|�4��=��5������YV�i{�J"���]�^�H�9��](�L�<O�C~�_<똠��c�;��E`Zx����ؠR���$���2�aqB�h�4-��V���+a��W���^U�vi��
y��ҿ�./ՎQd��/�u�7yF����J��
C���)q�N��s�b�N���a��Q�a 1�A9�oɹ��-��u�����nMn����G\��y�S�K?���,�9>���|��֦0PǛ$v̢��k)љ��"�4A'��?ʂ��+�,i�g������@Q[hijpJlR䊢��toT!���ܰ՟��l�����I�y5����KP!^v�%c&�GB�{���W�֠[p@p[�i.�_��2�^=#U��=NN��� 	��i�UM�#R�MK�4�X�T7^M��_�XT�'&���c���ajTM���.�Dg+^I��/1���gW��B7m�澡������#Y0��Z]�RdN��	}��#}�8�G<�/�2k�D��c��xkk���آ
��c4��
��@�y�:N�Ͳ���n\���X�#]�?�.ߺ�$+��P�8�i���gl����k�d����D7P�B."��?4�dq*�}�Y�kQ�l/����t�����pTP�ka���r��m����@��&g!8ڿs���� ������a����gױx�#��Q3�OG����p:%���7�] .c���%L��TT�CkF	��_��s�n�An�U`o|�� (����6	�� /� 7���+��,�es%�{z��t����GB�(�Z�Þ}(<v���*�i��LW�ʟV(Z�9�Y����g��X�Ѕͪ�򱟖A�C��d�_���o�H��P�[�B�������l��b�؄��KP�c��%��ߌ��Y��f��*%��}]�+DSZt�Ư��j�P_����,e&������͑�d.Z���j��Q�JX�Uk���!�ԥ�cuKi}����#�S�>�&�x��mH(^~�>LA ���N �$^�c���Ico��o���� }��(�� T&�����u���O��b�IC���|+j��k悸�KOAh���`�X ���^ͪd_]rT�,N��/�� U@
� �^��F->	1��p��n���)��n���Z��)D��e���}��
@���~���aTO��5ZA��L�J��}�ә~�t�V*�&��Ͼ$�9���3���5�n��W�&�R�;*������A�����v�D?Zn��c�eE�W�oi�B& �|͇8?��������g��)`�`�ҥ8�K7�]��E�:�}��B�p��8��`���i�ĥY*��n�V��Y)ݘ�@�	��_�x/�d��o���.5˃]O�������n���J�`]��ʌ͆�*-��:�HV�b����5\\� P+��M����#q�h|�����bR(BQ��V���8\�Ǌ��&bD�.���Zo�Tp$"�R�ޛ�f�d��8�?�˂rmw�h����IY��hg\�<E4���J�7�?�Ǥ������z�������C� "�+T�6�)$Jg_��Ϥ����j������V�5thx�U{��iT���JC��U!L��l`R���w��p���X�7�X���-Z	��X���k�=YS�K��a%�'�f�`�4�%�v�V�Tjg�j���,�,�������6�����
�� %A��O�ܾ�6�5h�&8-�Y��w�w�:��؋���bJa�g3�|�u��N�Yw��^��$�
�D��H����K�e4�o�����4Q@}q&�)G�&�x�����eUu�[��= �!�1�$c#x{�d�[��A�%Hr{.J��*S1 �J���T�`d�7�[��a�$yL���2�*Y�F��L2�k�yOk��Ŏ��݄�]/��dO�%;�q��q���9���b��b�H�����ns�)�U��1�f�N��1l!@���2�9@ۛH���%^�Sݏm���)Q,��D������	�	P;j�/��v_S(���ĤD����=�Z�B�yC���-���xݕB8C
��9������5��-d�%ԓ0b��yG�r����Ô�Ǚ��2��2Lv��n���/��?fb���=�
���ғŇ�a��_�x�����Bu�+���<w�Jl&���D�U�5�6y�\��uڄM>6��L�J�徾~J���J)ʏ�:�}ڿ��\������S�-gJ�|M�(�=�a��݃��[�l�&Z�+���-��B�I��C�.�ӵ�l_�S��#��i�-U�����V;�BW����]A��v�k���.�$��s�|�O��{��Пx9z����3r�Ǽ���9�����$CL���k�O�T-���\�a7ݴ�!�W�Tn�D���B+< ����Ҍ|�?,����N�1�ʦ���S�kb�pV8�z!��$�@��?�t�ɦ��CZ?�Z�%�G-�K�m�BƔ3��)�A�����%W��� �|z�ץkt~������8�~��M8�օE�+��V7��ScJ.���^Q㿲���l)t�g��u�X�$��^���@a���b��.¹�j ,e��)x�0#��(�#�!t�	#�s<6�X&�G�e�FtH+�K�����Eu��;���V�=��k�e�;���`�PB)]k�ݤC,�
�)?��9�"O����MQW�DmX}��y��/���E�0E	KՆ��Fx~�ς��Zd�.Lh��L�D����̹����A�v	y�����7v�-��X7i-��Ϯ\խ�[�:ur��X��g��-6����[��,��_����'�D	�<���h��)JI�.�vL~�3�w�>���"y����"ǘL��)N�wL{�����p��|J}��6L�!؂�7g��"G�VuC�=]��u$��>��lalU�/n��;_DHm�d��
n�K��sr]YJp���Tʽ!�l+d���N1��]Z�H�υ΁T���Y�� �-�H��\`:r�R:�_ٷo~�ȸ�B]�����ihgw.h��crǼ�Y^)�P2?�/�tu��Q!bO�[K�'��z��Y��]�i�['��R����G��^'u!��j� GKM���r����Q���:��	���u���X|���=g]�[?����4��w��[�x��4�^�k�����4ߩ�2Y��N�h� 1��S5L΄te%��ͫQ��B6�hi��/=��,_�V����"��&>�eavL�i=p{Rb����?1&յ��S=����j�C�����:>�P9s��3���C�_,E����r{5�������X�Ա�9T4���m���D��^P@�E+x�Lrp�M�!��� ξ¹��}���_��%2�(-5�q��Ua$�uW�`�������-.k�o�X��ui�A��n���_��p7�Џ�G��a}���o�998�C�x�ե|�TB��@���{�Ne�\�c8���٠�D<я�2��G�c�M�������;�_����|?+f6v���m����M�`�5��`�飽�T�u:��<oY�M�Tg�6��(̚5���_�"��Y��
B��uP���Ngs(�Ba�	�c�nߺ|L�[<�&Wh�U��ti�]K��(o��V���/����;�|,v;�k�zL�|�[t?`��I2�6��v��q�ϣ�%4��ma��1���$e�3Ho��\������rX�TG��br媃o9C��%s��8��� L���G���rUf�`C��a԰���Rʿ�ĵ���IN|z=��L�px�U���P����ʒN5��� ��[V6V �L�H���bA���M�D�i�q����b���F�U����Ƕå��g-n~A2u�bX!(��)���A���*��ݨ~#$4��x�f\��ؕ ��ʎ7��j!�Q�90�*"6�� <=�n���1�+���6?�6���%<�?E�g��n��p1���Q�I�?����e�Uӷ���ܔ�u?|�S<�rG��[��Ĵ���F�>7� �4��f����_���@Z��	���!�w��k��g�c�7^;����uU�4���&�9�F���O�<%�p���M�=h�^I�_b�^��u�$Sg�7I-�����.ė���Kp2cH�5;D�`K�^/l��0oM�ĕY{s��(颜p��,�J�a�:�Z;��
DV�G�3�o�u�����O�( �X֢>[f�I�Vazl�G���>bP!�
�O2������&�(���|�������tM�rѵc�q�n7@Q�t�(����ř���K.���c�iH
E��2��Df��d�m�ApsX��W�`_һ�6���W�S�y��;�ƅЙ%�U�,i��6�h��?g�y �o�v޶���(NG�bϞ~���WW���[��i����c)S�L�1�fEԴ�;_Q����c��[?<���f���f
�N���q[5$h��`��Hw�$n����Y�c��~�?py��+1�	�r�^�Y������0К��8���QX$��("���� ��`�l�M�3�r����w���b�!��}
<��ۑ��h�d��(-����4�14bnꆴΈm���/d+���8��[���FJ��U�����r-w[2��v�E̍H�%����N/8�������2�[1�[.��%a��FR,|�\�.���0 �I]�@W)�IF?�v�? �L=����U_���l��(�d!� LɄ����1��l�R���+�:���\�"�@�΋��NB��`À�"���j�/1'&ߕ5�GXA�"x\+������>��X:8��V�)U����w��*A�����1F�a���C#�����-�BU�(�,�{��c��Oy�u
y��O�f��	mp1!�Z]���EiC�]HkM�@�%���4�G��ZU]Yʙ��8�T�b ���cX�U���x�MH�Vw�c�쀎&��a0˖L��$_���,z��{k$�_̮2�b����p�5�Ҏ�E�+;p~�l����C����Frc��,��\��E�ʵ(D|����f�{��������>V��Ѝ_�����t�,&�7~C�Bӧ�Y,�uy�L�3�� �B/��ǘ���,B�r�w�V��.����&��8x���Y�e;����|Ԥ�Y��B��J�~=`b��,�-�G���րe��i�8�*�q�F�:`��a��+�1�D��z7��iN=F���;����#�\�#��3��ƕ���ݯ+a����gZl��n��Sd&g�W�Y�z�[ �� C,^��Ů����j�A�5�:]���m��f��V�}?P���'�:ENͦ�}{68��������V���t����b�����\���i��0�{� ��QŃY�����O��'�J�W�B}�~lg\�b����^�+�}=ѕ�b|S�V�2��jb��,w�8v����4� #��e�?����Yf�g��;5N�P�7�~u�@��/�f�\덚&�<_jQ�(����� //\_�:�`��,�(���4+�U�S�/��3���a����騻���
U{������z�,6dTr	u����g4���@ N_���R5#�
ĕ^`$�9�|�!�u�nT�5�[��t{�Jh��t��/�<����l��"���<�mX�q�R�KY?ys�$�	��[�I�r�;<��G����M�G9l>�K�}�����2�nt���zGH�  4[�F�@v؀k�=&�JjG	��I,����͟W�K��*�N�c���	�e��Ok��������oeN�'��oOj��W��^g#}����)g&���=B�0��`�!HΜ�2fX�m/�1x��j!qH|N)O�6�sh��}�t/4�")����n^k�kcMM!y��pw#�h��r��ju�dSI�6���)E��0��	�<�����u��>��.#��iҫY��v�[g�����=�P-�b�[&l�����|y$���m��:d紫�ScV�r�9���̕��@.�>D��`ǎ�G"�W<�q�g[_	�ǀ B|�����k�[@�lEі�QY��.����ɒ~�-�ĥ��WW���\�$jyIY�B.���e�R\�g��D.D&��� k�Q��Ѫ�������	��H��C\���Ez���Z
�P,8�����'D80 �0����vv������{ߧ�V�	|�fyl �"k��t�\������֘��GS��(q�/�HQ+�Wa�-��*�;��3I��߶E�� ˘���x>��W}�~�9D�+�-�k��:��ȰwF}���v�N-����%;J��M^푙^	��t��� 3jl��1İf�9�����#K�q|��D�On��ѡ~��2���'Lx�Z/&׉�6[��_<��&_�1��������������}�#��ח�27�������"����Ԅ���E��1h�D	����R��<����.�9=�pm��S�L��r�d,:� '��C�g{ơ	ϼ%��xPD��m��ôt-/dc�VT�~Lj�_��U�?�{_oZ`?���qJ��(If<���;�^�JM:�%�������U��`H΃艳g��P3{t��[�Z����j<*^K���]}�%�u�S���ZN>&��p�����h�[��":��e�sA��[����]�<�&N�2=�4�3u:�P��i�4��ކ��Ld��ۢ93_������_�> @�3��AA�g����^����⯃��. C<��BE�b9�$��0�:^�&�сAa��*�j[����,�/h;I\Dg�,BMMr��r������!M�]���n�q��j�Rf&F���'���$Ã:����+jq�"F��<�-Uq<:����̪�\L��3A���v���AF"�5t��k��p�my���E���	 &I�y��/��k�����HSS�OeaB0>�����4� �Ó���e�����sOF숶J������b�a.�Z��H�K�#[z�-�5��o@���=�zm%�l>k�筳�;3����E@�U]pS��� ������(���]�K�L�π�,?q��@��hեS�;f��!y�$���|�kG<�����V�?��U����|iV�gE�L5�гa#AQ�E�~ZD1���B��$�!(w��6)Z=/��\���5U�{3�)�ل���,��>)��k���{
88��	��n �y�2�,��H{��FV��C���zc�U�`�/@�/�m,�`��O���W���(��������B��EQҖ�@�n�C04,��$<��{���!LNٻ�k�u�5tA�<�,|�Z�C�]��Q�a*���EdO�C[ݖ�K���/+���5f̞U�-�R���s��X+|�u�6A-����a�ei���(���o:�Q��"4M�H�X�̘�G-� �e�M��yC�ն�d��^g![���VNj~����\>�O���V����n��
�
OG��Ϙ��\R��7
���k�Zv^��eq~$�GtR�A%����}XR�K`'y�'Y�H_�ɮ��1a��̺+"7��.�(A1�_� �J�]�ob�2y�y�/Wd���F�G=��O�"ܐ�1�Smb.D�l
y��SRd�t����dY�܈�	}�p������&\���v﨟ntYY!�e�I�~�f���y�\sU~\��/c<��b̓�D�q^:��G�Y���N��kU�y�'Y�Ȉ�k�w����4-�2le�g:�9$� �t��%)���*��}�/`�t	��~�k����o��q��3%'��P�^��,R�$�nQ��[8���F1o�z�)]��ˬ���/�L�8�z��`�F��������8�j(q[\����vt��rC��#~�$�����Gg�n:�8&w6�4����s�~��D}�tk�ʁ������̸�?)M#�;�Ӑ;��Ӗ�,.5?�C��4,���������Q��}���l����{��R3�z,}�[[c~���X&aߢ2�7�"�A����g#�����{��$���J?@=�8yQ��x�8��^p85�k�|/PגR2:�W ɉK��|#�����i��H}�؆�J8��xpm��&�7X�ɩ�t&;��RۿżEޏ-e8��h����J���B�p�ӫR}��B���ק\(��F�/�^�z��ݶE%�i���>Dqh0�5[�(�����F:
�Pd�W<��	��`����#.�=����}���=��ae*|b@�i�Z����K� k߉��K3]��!��H�ﲫ�}�/C}�C���{�hpWq�%%�G�6�B���b�'sǁ��S*:��%��*r{��V
�-���7B����2���OH���i|^��9�I�7멷��X��"@����K}�xtj/��c��R�f8�&�o$jXJwqM?�_���)��Ns`�A	
s�O��iG$�-+��uo���I��{H�����c�m��%\�/A�n���ʞ=_����{��Z|�ZN���ϳ�cX��%�>;V!a�	*�9�őyC�_~�s���I�!��˵��m�ܘw!4�����u%m˹���S�\<���:5����
�L�)|-�9��8迣m��W����������%W%r��II_8�/l�ǳ§��}�C�Bv=*ɨ!�74�����������!����=�<K�&�N����[���3v�����Ǯ���s�%��]8����s��t'�ѕ��g1+w�ă�[��dwX�p"9+��!��H��0(�U4���Vd�BJt��=)N+����q#���//<h@�B�(	 lt�� 1�r��(qy]��?i�Z�@a Ǚ�`�c�c���"iP��n=�4�ǩXV"�J?�̽�ɋt��!0�Q|SV�� ���=��[��0�$��묋\��̐��qqd��/orӮ]�W��3[���M��O"5n\��,9uA�,0 >���2��%3X�/þ}�YH��^
3*��4vkĐ�;ꀤG`�m���[�TnS��pi�wP#�܍<��/��/QY���. 6L��z�Xo�+���"Y������ʅ��ٝ�q�0:f WDi�r�D(l���* s�ۏͳ�Tk�:��*����B@^�y�`�N���X<th�2���"���������ς@H&E�*��'I�fq����X�D\�w#I��<�㳙�d�V�9kܘv��O&�.� ��@�,��qF=�X�M��J���=�0���@)�1Q�~o"RP��F~���K����f(�x;� {JT�J)]�M��i����:K�c�[w�籲�����k����F�.%̜�+D�\�}�<�2��σ��uzЏw�\W,��s;n�R6!y�smc�A^��&����^�=r�qR�)b�c�M�;B�8��I�3�{�{