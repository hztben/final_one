  --Example instantiation for system 'nios2'
  nios2_inst : nios2
    port map(
      address_to_the_cfi_flash_0 => address_to_the_cfi_flash_0,
      data_to_and_from_the_cfi_flash_0 => data_to_and_from_the_cfi_flash_0,
      dclk_from_the_epcs_flash_controller_0 => dclk_from_the_epcs_flash_controller_0,
      out_port_from_the_addr => out_port_from_the_addr,
      out_port_from_the_addr2 => out_port_from_the_addr2,
      out_port_from_the_addr3 => out_port_from_the_addr3,
      out_port_from_the_addr4 => out_port_from_the_addr4,
      out_port_from_the_pio_1 => out_port_from_the_pio_1,
      out_port_from_the_pio_2 => out_port_from_the_pio_2,
      out_port_from_the_pio_3 => out_port_from_the_pio_3,
      out_port_from_the_pio_4 => out_port_from_the_pio_4,
      out_port_from_the_wr => out_port_from_the_wr,
      out_port_from_the_wr2 => out_port_from_the_wr2,
      out_port_from_the_wr3 => out_port_from_the_wr3,
      out_port_from_the_wr4 => out_port_from_the_wr4,
      read_n_to_the_cfi_flash_0 => read_n_to_the_cfi_flash_0,
      sce_from_the_epcs_flash_controller_0 => sce_from_the_epcs_flash_controller_0,
      scl_pad_io_to_and_from_the_opencores_i2c_fbm320 => scl_pad_io_to_and_from_the_opencores_i2c_fbm320,
      scl_pad_io_to_and_from_the_opencores_i2c_jy901 => scl_pad_io_to_and_from_the_opencores_i2c_jy901,
      sda_pad_io_to_and_from_the_opencores_i2c_fbm320 => sda_pad_io_to_and_from_the_opencores_i2c_fbm320,
      sda_pad_io_to_and_from_the_opencores_i2c_jy901 => sda_pad_io_to_and_from_the_opencores_i2c_jy901,
      sdo_from_the_epcs_flash_controller_0 => sdo_from_the_epcs_flash_controller_0,
      select_n_to_the_cfi_flash_0 => select_n_to_the_cfi_flash_0,
      txd_from_the_HC_12 => txd_from_the_HC_12,
      txd_from_the_US_100_UART => txd_from_the_US_100_UART,
      write_n_to_the_cfi_flash_0 => write_n_to_the_cfi_flash_0,
      zs_addr_from_the_sdram_0 => zs_addr_from_the_sdram_0,
      zs_ba_from_the_sdram_0 => zs_ba_from_the_sdram_0,
      zs_cas_n_from_the_sdram_0 => zs_cas_n_from_the_sdram_0,
      zs_cke_from_the_sdram_0 => zs_cke_from_the_sdram_0,
      zs_cs_n_from_the_sdram_0 => zs_cs_n_from_the_sdram_0,
      zs_dq_to_and_from_the_sdram_0 => zs_dq_to_and_from_the_sdram_0,
      zs_dqm_from_the_sdram_0 => zs_dqm_from_the_sdram_0,
      zs_ras_n_from_the_sdram_0 => zs_ras_n_from_the_sdram_0,
      zs_we_n_from_the_sdram_0 => zs_we_n_from_the_sdram_0,
      clk_0 => clk_0,
      data0_to_the_epcs_flash_controller_0 => data0_to_the_epcs_flash_controller_0,
      in_port_to_the_pio_0 => in_port_to_the_pio_0,
      reset_n => reset_n,
      rxd_to_the_HC_12 => rxd_to_the_HC_12,
      rxd_to_the_US_100_UART => rxd_to_the_US_100_UART
    );


